-- Copyright (C) 2022  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- ***************************************************************************
-- This file contains a Vhdl test bench template that is freely editable to   
-- suit user's needs .Comments are provided in each section to help the user  
-- fill out necessary details.                                                
-- ***************************************************************************
-- Generated on "03/14/2025 11:37:18"
                                                            
-- Vhdl Test Bench template for design  :  universal_register
-- 
-- Simulation tool : Questa Intel FPGA (VHDL)
-- 

LIBRARY ieee;                                               
USE ieee.std_logic_1164.all;                                

ENTITY tb_shift_register_universal8_prof IS
END tb_shift_register_universal8_prof;

ARCHITECTURE universal_register_arch OF tb_shift_register_universal8_prof IS
-- constants                                                 
-- signals                                                   
SIGNAL CLK : STD_LOGIC;
SIGNAL RSTn : STD_LOGIC;
SIGNAL SETn : STD_LOGIC;
SIGNAL SEL : STD_LOGIC_VECTOR(2 downto 0);
SIGNAL SSR : STD_LOGIC;
SIGNAL SSL : STD_LOGIC;
SIGNAL Pi : STD_LOGIC_VECTOR(7 downto 0);
SIGNAL Qo : STD_LOGIC_VECTOR(7 downto 0);
SIGNAL SOR : STD_LOGIC;
SIGNAL SOL : STD_LOGIC;

BEGIN
	UUT : entity work.shift_register_universal8
	PORT MAP (
-- list connections between master ports and signals
	CLK => CLK,
	RSTn => RSTn,
	SETn => SETn,
    SEL => SEL,
    SSR => SSR,
    SSL => SSL,
    Pi => Pi,
    Qo => Qo,
    SOR => SOR,
    SOL => SOL
	);

stimuli : process
    begin
    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1/2803" severity error;
    assert SOR = '0' report "Error in test case #1/2803" severity error;
    assert SOL = '0' report "Error in test case #1/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2/2803" severity error;
    assert SOR = '0' report "Error in test case #2/2803" severity error;
    assert SOL = '0' report "Error in test case #2/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #3/2803" severity error;
    assert SOR = '0' report "Error in test case #3/2803" severity error;
    assert SOL = '0' report "Error in test case #3/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #4/2803" severity error;
    assert SOR = '0' report "Error in test case #4/2803" severity error;
    assert SOL = '0' report "Error in test case #4/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #5/2803" severity error;
    assert SOR = '0' report "Error in test case #5/2803" severity error;
    assert SOL = '0' report "Error in test case #5/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #6/2803" severity error;
    assert SOR = '0' report "Error in test case #6/2803" severity error;
    assert SOL = '0' report "Error in test case #6/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #7/2803" severity error;
    assert SOR = '0' report "Error in test case #7/2803" severity error;
    assert SOL = '0' report "Error in test case #7/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #8/2803" severity error;
    assert SOR = '0' report "Error in test case #8/2803" severity error;
    assert SOL = '0' report "Error in test case #8/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #9/2803" severity error;
    assert SOR = '0' report "Error in test case #9/2803" severity error;
    assert SOL = '0' report "Error in test case #9/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #10/2803" severity error;
    assert SOR = '0' report "Error in test case #10/2803" severity error;
    assert SOL = '0' report "Error in test case #10/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #11/2803" severity error;
    assert SOR = '0' report "Error in test case #11/2803" severity error;
    assert SOL = '0' report "Error in test case #11/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #12/2803" severity error;
    assert SOR = '0' report "Error in test case #12/2803" severity error;
    assert SOL = '0' report "Error in test case #12/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #13/2803" severity error;
    assert SOR = '0' report "Error in test case #13/2803" severity error;
    assert SOL = '0' report "Error in test case #13/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #14/2803" severity error;
    assert SOR = '0' report "Error in test case #14/2803" severity error;
    assert SOL = '0' report "Error in test case #14/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #15/2803" severity error;
    assert SOR = '0' report "Error in test case #15/2803" severity error;
    assert SOL = '0' report "Error in test case #15/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #16/2803" severity error;
    assert SOR = '0' report "Error in test case #16/2803" severity error;
    assert SOL = '0' report "Error in test case #16/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #17/2803" severity error;
    assert SOR = '0' report "Error in test case #17/2803" severity error;
    assert SOL = '0' report "Error in test case #17/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #18/2803" severity error;
    assert SOR = '0' report "Error in test case #18/2803" severity error;
    assert SOL = '0' report "Error in test case #18/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #19/2803" severity error;
    assert SOR = '0' report "Error in test case #19/2803" severity error;
    assert SOL = '0' report "Error in test case #19/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #20/2803" severity error;
    assert SOR = '0' report "Error in test case #20/2803" severity error;
    assert SOL = '0' report "Error in test case #20/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #21/2803" severity error;
    assert SOR = '0' report "Error in test case #21/2803" severity error;
    assert SOL = '0' report "Error in test case #21/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #22/2803" severity error;
    assert SOR = '0' report "Error in test case #22/2803" severity error;
    assert SOL = '0' report "Error in test case #22/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #23/2803" severity error;
    assert SOR = '0' report "Error in test case #23/2803" severity error;
    assert SOL = '0' report "Error in test case #23/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #24/2803" severity error;
    assert SOR = '0' report "Error in test case #24/2803" severity error;
    assert SOL = '0' report "Error in test case #24/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #25/2803" severity error;
    assert SOR = '0' report "Error in test case #25/2803" severity error;
    assert SOL = '0' report "Error in test case #25/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #26/2803" severity error;
    assert SOR = '0' report "Error in test case #26/2803" severity error;
    assert SOL = '0' report "Error in test case #26/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #27/2803" severity error;
    assert SOR = '0' report "Error in test case #27/2803" severity error;
    assert SOL = '0' report "Error in test case #27/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #28/2803" severity error;
    assert SOR = '0' report "Error in test case #28/2803" severity error;
    assert SOL = '0' report "Error in test case #28/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #29/2803" severity error;
    assert SOR = '0' report "Error in test case #29/2803" severity error;
    assert SOL = '0' report "Error in test case #29/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #30/2803" severity error;
    assert SOR = '0' report "Error in test case #30/2803" severity error;
    assert SOL = '0' report "Error in test case #30/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #31/2803" severity error;
    assert SOR = '0' report "Error in test case #31/2803" severity error;
    assert SOL = '0' report "Error in test case #31/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #32/2803" severity error;
    assert SOR = '0' report "Error in test case #32/2803" severity error;
    assert SOL = '0' report "Error in test case #32/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #33/2803" severity error;
    assert SOR = '0' report "Error in test case #33/2803" severity error;
    assert SOL = '0' report "Error in test case #33/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #34/2803" severity error;
    assert SOR = '0' report "Error in test case #34/2803" severity error;
    assert SOL = '0' report "Error in test case #34/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #35/2803" severity error;
    assert SOR = '0' report "Error in test case #35/2803" severity error;
    assert SOL = '0' report "Error in test case #35/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #36/2803" severity error;
    assert SOR = '0' report "Error in test case #36/2803" severity error;
    assert SOL = '0' report "Error in test case #36/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #37/2803" severity error;
    assert SOR = '0' report "Error in test case #37/2803" severity error;
    assert SOL = '0' report "Error in test case #37/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #38/2803" severity error;
    assert SOR = '0' report "Error in test case #38/2803" severity error;
    assert SOL = '0' report "Error in test case #38/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #39/2803" severity error;
    assert SOR = '0' report "Error in test case #39/2803" severity error;
    assert SOL = '0' report "Error in test case #39/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #40/2803" severity error;
    assert SOR = '0' report "Error in test case #40/2803" severity error;
    assert SOL = '0' report "Error in test case #40/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #41/2803" severity error;
    assert SOR = '0' report "Error in test case #41/2803" severity error;
    assert SOL = '0' report "Error in test case #41/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #42/2803" severity error;
    assert SOR = '0' report "Error in test case #42/2803" severity error;
    assert SOL = '0' report "Error in test case #42/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #43/2803" severity error;
    assert SOR = '0' report "Error in test case #43/2803" severity error;
    assert SOL = '0' report "Error in test case #43/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #44/2803" severity error;
    assert SOR = '0' report "Error in test case #44/2803" severity error;
    assert SOL = '0' report "Error in test case #44/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #45/2803" severity error;
    assert SOR = '0' report "Error in test case #45/2803" severity error;
    assert SOL = '0' report "Error in test case #45/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #46/2803" severity error;
    assert SOR = '0' report "Error in test case #46/2803" severity error;
    assert SOL = '0' report "Error in test case #46/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #47/2803" severity error;
    assert SOR = '0' report "Error in test case #47/2803" severity error;
    assert SOL = '0' report "Error in test case #47/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #48/2803" severity error;
    assert SOR = '0' report "Error in test case #48/2803" severity error;
    assert SOL = '0' report "Error in test case #48/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #49/2803" severity error;
    assert SOR = '0' report "Error in test case #49/2803" severity error;
    assert SOL = '0' report "Error in test case #49/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #50/2803" severity error;
    assert SOR = '0' report "Error in test case #50/2803" severity error;
    assert SOL = '0' report "Error in test case #50/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #51/2803" severity error;
    assert SOR = '0' report "Error in test case #51/2803" severity error;
    assert SOL = '0' report "Error in test case #51/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #52/2803" severity error;
    assert SOR = '0' report "Error in test case #52/2803" severity error;
    assert SOL = '0' report "Error in test case #52/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #53/2803" severity error;
    assert SOR = '0' report "Error in test case #53/2803" severity error;
    assert SOL = '0' report "Error in test case #53/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #54/2803" severity error;
    assert SOR = '0' report "Error in test case #54/2803" severity error;
    assert SOL = '0' report "Error in test case #54/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #55/2803" severity error;
    assert SOR = '0' report "Error in test case #55/2803" severity error;
    assert SOL = '0' report "Error in test case #55/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #56/2803" severity error;
    assert SOR = '0' report "Error in test case #56/2803" severity error;
    assert SOL = '0' report "Error in test case #56/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #57/2803" severity error;
    assert SOR = '0' report "Error in test case #57/2803" severity error;
    assert SOL = '0' report "Error in test case #57/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #58/2803" severity error;
    assert SOR = '0' report "Error in test case #58/2803" severity error;
    assert SOL = '0' report "Error in test case #58/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #59/2803" severity error;
    assert SOR = '0' report "Error in test case #59/2803" severity error;
    assert SOL = '0' report "Error in test case #59/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #60/2803" severity error;
    assert SOR = '0' report "Error in test case #60/2803" severity error;
    assert SOL = '0' report "Error in test case #60/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #61/2803" severity error;
    assert SOR = '0' report "Error in test case #61/2803" severity error;
    assert SOL = '0' report "Error in test case #61/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #62/2803" severity error;
    assert SOR = '0' report "Error in test case #62/2803" severity error;
    assert SOL = '0' report "Error in test case #62/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #63/2803" severity error;
    assert SOR = '0' report "Error in test case #63/2803" severity error;
    assert SOL = '0' report "Error in test case #63/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #64/2803" severity error;
    assert SOR = '0' report "Error in test case #64/2803" severity error;
    assert SOL = '0' report "Error in test case #64/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #65/2803" severity error;
    assert SOR = '0' report "Error in test case #65/2803" severity error;
    assert SOL = '0' report "Error in test case #65/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #66/2803" severity error;
    assert SOR = '0' report "Error in test case #66/2803" severity error;
    assert SOL = '0' report "Error in test case #66/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #67/2803" severity error;
    assert SOR = '0' report "Error in test case #67/2803" severity error;
    assert SOL = '0' report "Error in test case #67/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #68/2803" severity error;
    assert SOR = '0' report "Error in test case #68/2803" severity error;
    assert SOL = '0' report "Error in test case #68/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #69/2803" severity error;
    assert SOR = '0' report "Error in test case #69/2803" severity error;
    assert SOL = '0' report "Error in test case #69/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #70/2803" severity error;
    assert SOR = '0' report "Error in test case #70/2803" severity error;
    assert SOL = '0' report "Error in test case #70/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #71/2803" severity error;
    assert SOR = '0' report "Error in test case #71/2803" severity error;
    assert SOL = '0' report "Error in test case #71/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #72/2803" severity error;
    assert SOR = '0' report "Error in test case #72/2803" severity error;
    assert SOL = '0' report "Error in test case #72/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #73/2803" severity error;
    assert SOR = '0' report "Error in test case #73/2803" severity error;
    assert SOL = '0' report "Error in test case #73/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #74/2803" severity error;
    assert SOR = '0' report "Error in test case #74/2803" severity error;
    assert SOL = '0' report "Error in test case #74/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #75/2803" severity error;
    assert SOR = '0' report "Error in test case #75/2803" severity error;
    assert SOL = '0' report "Error in test case #75/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #76/2803" severity error;
    assert SOR = '0' report "Error in test case #76/2803" severity error;
    assert SOL = '0' report "Error in test case #76/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #77/2803" severity error;
    assert SOR = '0' report "Error in test case #77/2803" severity error;
    assert SOL = '0' report "Error in test case #77/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #78/2803" severity error;
    assert SOR = '0' report "Error in test case #78/2803" severity error;
    assert SOL = '0' report "Error in test case #78/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #79/2803" severity error;
    assert SOR = '0' report "Error in test case #79/2803" severity error;
    assert SOL = '0' report "Error in test case #79/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #80/2803" severity error;
    assert SOR = '0' report "Error in test case #80/2803" severity error;
    assert SOL = '0' report "Error in test case #80/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #81/2803" severity error;
    assert SOR = '0' report "Error in test case #81/2803" severity error;
    assert SOL = '0' report "Error in test case #81/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #82/2803" severity error;
    assert SOR = '0' report "Error in test case #82/2803" severity error;
    assert SOL = '0' report "Error in test case #82/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #83/2803" severity error;
    assert SOR = '0' report "Error in test case #83/2803" severity error;
    assert SOL = '0' report "Error in test case #83/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #84/2803" severity error;
    assert SOR = '0' report "Error in test case #84/2803" severity error;
    assert SOL = '0' report "Error in test case #84/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #85/2803" severity error;
    assert SOR = '0' report "Error in test case #85/2803" severity error;
    assert SOL = '0' report "Error in test case #85/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #86/2803" severity error;
    assert SOR = '0' report "Error in test case #86/2803" severity error;
    assert SOL = '0' report "Error in test case #86/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #87/2803" severity error;
    assert SOR = '0' report "Error in test case #87/2803" severity error;
    assert SOL = '0' report "Error in test case #87/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #88/2803" severity error;
    assert SOR = '0' report "Error in test case #88/2803" severity error;
    assert SOL = '0' report "Error in test case #88/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #89/2803" severity error;
    assert SOR = '0' report "Error in test case #89/2803" severity error;
    assert SOL = '0' report "Error in test case #89/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #90/2803" severity error;
    assert SOR = '0' report "Error in test case #90/2803" severity error;
    assert SOL = '0' report "Error in test case #90/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #91/2803" severity error;
    assert SOR = '0' report "Error in test case #91/2803" severity error;
    assert SOL = '0' report "Error in test case #91/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #92/2803" severity error;
    assert SOR = '0' report "Error in test case #92/2803" severity error;
    assert SOL = '0' report "Error in test case #92/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #93/2803" severity error;
    assert SOR = '0' report "Error in test case #93/2803" severity error;
    assert SOL = '0' report "Error in test case #93/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #94/2803" severity error;
    assert SOR = '0' report "Error in test case #94/2803" severity error;
    assert SOL = '0' report "Error in test case #94/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #95/2803" severity error;
    assert SOR = '0' report "Error in test case #95/2803" severity error;
    assert SOL = '0' report "Error in test case #95/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #96/2803" severity error;
    assert SOR = '0' report "Error in test case #96/2803" severity error;
    assert SOL = '0' report "Error in test case #96/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #97/2803" severity error;
    assert SOR = '0' report "Error in test case #97/2803" severity error;
    assert SOL = '0' report "Error in test case #97/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #98/2803" severity error;
    assert SOR = '0' report "Error in test case #98/2803" severity error;
    assert SOL = '0' report "Error in test case #98/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #99/2803" severity error;
    assert SOR = '0' report "Error in test case #99/2803" severity error;
    assert SOL = '0' report "Error in test case #99/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #100/2803" severity error;
    assert SOR = '0' report "Error in test case #100/2803" severity error;
    assert SOL = '0' report "Error in test case #100/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #101/2803" severity error;
    assert SOR = '0' report "Error in test case #101/2803" severity error;
    assert SOL = '0' report "Error in test case #101/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #102/2803" severity error;
    assert SOR = '0' report "Error in test case #102/2803" severity error;
    assert SOL = '0' report "Error in test case #102/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #103/2803" severity error;
    assert SOR = '0' report "Error in test case #103/2803" severity error;
    assert SOL = '0' report "Error in test case #103/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #104/2803" severity error;
    assert SOR = '0' report "Error in test case #104/2803" severity error;
    assert SOL = '0' report "Error in test case #104/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #105/2803" severity error;
    assert SOR = '0' report "Error in test case #105/2803" severity error;
    assert SOL = '0' report "Error in test case #105/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #106/2803" severity error;
    assert SOR = '0' report "Error in test case #106/2803" severity error;
    assert SOL = '0' report "Error in test case #106/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #107/2803" severity error;
    assert SOR = '0' report "Error in test case #107/2803" severity error;
    assert SOL = '0' report "Error in test case #107/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #108/2803" severity error;
    assert SOR = '0' report "Error in test case #108/2803" severity error;
    assert SOL = '0' report "Error in test case #108/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #109/2803" severity error;
    assert SOR = '0' report "Error in test case #109/2803" severity error;
    assert SOL = '0' report "Error in test case #109/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #110/2803" severity error;
    assert SOR = '0' report "Error in test case #110/2803" severity error;
    assert SOL = '0' report "Error in test case #110/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #111/2803" severity error;
    assert SOR = '0' report "Error in test case #111/2803" severity error;
    assert SOL = '0' report "Error in test case #111/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #112/2803" severity error;
    assert SOR = '0' report "Error in test case #112/2803" severity error;
    assert SOL = '0' report "Error in test case #112/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #113/2803" severity error;
    assert SOR = '0' report "Error in test case #113/2803" severity error;
    assert SOL = '0' report "Error in test case #113/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #114/2803" severity error;
    assert SOR = '0' report "Error in test case #114/2803" severity error;
    assert SOL = '0' report "Error in test case #114/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #115/2803" severity error;
    assert SOR = '0' report "Error in test case #115/2803" severity error;
    assert SOL = '0' report "Error in test case #115/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #116/2803" severity error;
    assert SOR = '0' report "Error in test case #116/2803" severity error;
    assert SOL = '0' report "Error in test case #116/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #117/2803" severity error;
    assert SOR = '0' report "Error in test case #117/2803" severity error;
    assert SOL = '0' report "Error in test case #117/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #118/2803" severity error;
    assert SOR = '0' report "Error in test case #118/2803" severity error;
    assert SOL = '0' report "Error in test case #118/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #119/2803" severity error;
    assert SOR = '0' report "Error in test case #119/2803" severity error;
    assert SOL = '0' report "Error in test case #119/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #120/2803" severity error;
    assert SOR = '0' report "Error in test case #120/2803" severity error;
    assert SOL = '0' report "Error in test case #120/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #121/2803" severity error;
    assert SOR = '0' report "Error in test case #121/2803" severity error;
    assert SOL = '0' report "Error in test case #121/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #122/2803" severity error;
    assert SOR = '0' report "Error in test case #122/2803" severity error;
    assert SOL = '0' report "Error in test case #122/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #123/2803" severity error;
    assert SOR = '0' report "Error in test case #123/2803" severity error;
    assert SOL = '0' report "Error in test case #123/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #124/2803" severity error;
    assert SOR = '0' report "Error in test case #124/2803" severity error;
    assert SOL = '0' report "Error in test case #124/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #125/2803" severity error;
    assert SOR = '0' report "Error in test case #125/2803" severity error;
    assert SOL = '0' report "Error in test case #125/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #126/2803" severity error;
    assert SOR = '0' report "Error in test case #126/2803" severity error;
    assert SOL = '0' report "Error in test case #126/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #127/2803" severity error;
    assert SOR = '0' report "Error in test case #127/2803" severity error;
    assert SOL = '0' report "Error in test case #127/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #128/2803" severity error;
    assert SOR = '0' report "Error in test case #128/2803" severity error;
    assert SOL = '0' report "Error in test case #128/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #129/2803" severity error;
    assert SOR = '0' report "Error in test case #129/2803" severity error;
    assert SOL = '0' report "Error in test case #129/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #130/2803" severity error;
    assert SOR = '0' report "Error in test case #130/2803" severity error;
    assert SOL = '0' report "Error in test case #130/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #131/2803" severity error;
    assert SOR = '0' report "Error in test case #131/2803" severity error;
    assert SOL = '0' report "Error in test case #131/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #132/2803" severity error;
    assert SOR = '0' report "Error in test case #132/2803" severity error;
    assert SOL = '0' report "Error in test case #132/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #133/2803" severity error;
    assert SOR = '0' report "Error in test case #133/2803" severity error;
    assert SOL = '0' report "Error in test case #133/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #134/2803" severity error;
    assert SOR = '0' report "Error in test case #134/2803" severity error;
    assert SOL = '0' report "Error in test case #134/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #135/2803" severity error;
    assert SOR = '0' report "Error in test case #135/2803" severity error;
    assert SOL = '0' report "Error in test case #135/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #136/2803" severity error;
    assert SOR = '0' report "Error in test case #136/2803" severity error;
    assert SOL = '0' report "Error in test case #136/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #137/2803" severity error;
    assert SOR = '0' report "Error in test case #137/2803" severity error;
    assert SOL = '0' report "Error in test case #137/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #138/2803" severity error;
    assert SOR = '0' report "Error in test case #138/2803" severity error;
    assert SOL = '0' report "Error in test case #138/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #139/2803" severity error;
    assert SOR = '0' report "Error in test case #139/2803" severity error;
    assert SOL = '0' report "Error in test case #139/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #140/2803" severity error;
    assert SOR = '0' report "Error in test case #140/2803" severity error;
    assert SOL = '0' report "Error in test case #140/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #141/2803" severity error;
    assert SOR = '0' report "Error in test case #141/2803" severity error;
    assert SOL = '0' report "Error in test case #141/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #142/2803" severity error;
    assert SOR = '0' report "Error in test case #142/2803" severity error;
    assert SOL = '0' report "Error in test case #142/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #143/2803" severity error;
    assert SOR = '0' report "Error in test case #143/2803" severity error;
    assert SOL = '0' report "Error in test case #143/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #144/2803" severity error;
    assert SOR = '0' report "Error in test case #144/2803" severity error;
    assert SOL = '0' report "Error in test case #144/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #145/2803" severity error;
    assert SOR = '0' report "Error in test case #145/2803" severity error;
    assert SOL = '0' report "Error in test case #145/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #146/2803" severity error;
    assert SOR = '0' report "Error in test case #146/2803" severity error;
    assert SOL = '0' report "Error in test case #146/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #147/2803" severity error;
    assert SOR = '0' report "Error in test case #147/2803" severity error;
    assert SOL = '0' report "Error in test case #147/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #148/2803" severity error;
    assert SOR = '0' report "Error in test case #148/2803" severity error;
    assert SOL = '0' report "Error in test case #148/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #149/2803" severity error;
    assert SOR = '0' report "Error in test case #149/2803" severity error;
    assert SOL = '0' report "Error in test case #149/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #150/2803" severity error;
    assert SOR = '0' report "Error in test case #150/2803" severity error;
    assert SOL = '0' report "Error in test case #150/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #151/2803" severity error;
    assert SOR = '0' report "Error in test case #151/2803" severity error;
    assert SOL = '0' report "Error in test case #151/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #152/2803" severity error;
    assert SOR = '0' report "Error in test case #152/2803" severity error;
    assert SOL = '0' report "Error in test case #152/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #153/2803" severity error;
    assert SOR = '0' report "Error in test case #153/2803" severity error;
    assert SOL = '0' report "Error in test case #153/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #154/2803" severity error;
    assert SOR = '0' report "Error in test case #154/2803" severity error;
    assert SOL = '0' report "Error in test case #154/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #155/2803" severity error;
    assert SOR = '0' report "Error in test case #155/2803" severity error;
    assert SOL = '0' report "Error in test case #155/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #156/2803" severity error;
    assert SOR = '0' report "Error in test case #156/2803" severity error;
    assert SOL = '0' report "Error in test case #156/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #157/2803" severity error;
    assert SOR = '0' report "Error in test case #157/2803" severity error;
    assert SOL = '0' report "Error in test case #157/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #158/2803" severity error;
    assert SOR = '0' report "Error in test case #158/2803" severity error;
    assert SOL = '0' report "Error in test case #158/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #159/2803" severity error;
    assert SOR = '0' report "Error in test case #159/2803" severity error;
    assert SOL = '0' report "Error in test case #159/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #160/2803" severity error;
    assert SOR = '0' report "Error in test case #160/2803" severity error;
    assert SOL = '0' report "Error in test case #160/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #161/2803" severity error;
    assert SOR = '0' report "Error in test case #161/2803" severity error;
    assert SOL = '0' report "Error in test case #161/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #162/2803" severity error;
    assert SOR = '0' report "Error in test case #162/2803" severity error;
    assert SOL = '0' report "Error in test case #162/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #163/2803" severity error;
    assert SOR = '0' report "Error in test case #163/2803" severity error;
    assert SOL = '0' report "Error in test case #163/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #164/2803" severity error;
    assert SOR = '0' report "Error in test case #164/2803" severity error;
    assert SOL = '0' report "Error in test case #164/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #165/2803" severity error;
    assert SOR = '0' report "Error in test case #165/2803" severity error;
    assert SOL = '0' report "Error in test case #165/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #166/2803" severity error;
    assert SOR = '0' report "Error in test case #166/2803" severity error;
    assert SOL = '0' report "Error in test case #166/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #167/2803" severity error;
    assert SOR = '0' report "Error in test case #167/2803" severity error;
    assert SOL = '0' report "Error in test case #167/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #168/2803" severity error;
    assert SOR = '0' report "Error in test case #168/2803" severity error;
    assert SOL = '0' report "Error in test case #168/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #169/2803" severity error;
    assert SOR = '0' report "Error in test case #169/2803" severity error;
    assert SOL = '0' report "Error in test case #169/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #170/2803" severity error;
    assert SOR = '0' report "Error in test case #170/2803" severity error;
    assert SOL = '0' report "Error in test case #170/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #171/2803" severity error;
    assert SOR = '0' report "Error in test case #171/2803" severity error;
    assert SOL = '0' report "Error in test case #171/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #172/2803" severity error;
    assert SOR = '0' report "Error in test case #172/2803" severity error;
    assert SOL = '0' report "Error in test case #172/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #173/2803" severity error;
    assert SOR = '0' report "Error in test case #173/2803" severity error;
    assert SOL = '0' report "Error in test case #173/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #174/2803" severity error;
    assert SOR = '0' report "Error in test case #174/2803" severity error;
    assert SOL = '0' report "Error in test case #174/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #175/2803" severity error;
    assert SOR = '0' report "Error in test case #175/2803" severity error;
    assert SOL = '0' report "Error in test case #175/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #176/2803" severity error;
    assert SOR = '0' report "Error in test case #176/2803" severity error;
    assert SOL = '0' report "Error in test case #176/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #177/2803" severity error;
    assert SOR = '0' report "Error in test case #177/2803" severity error;
    assert SOL = '0' report "Error in test case #177/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #178/2803" severity error;
    assert SOR = '0' report "Error in test case #178/2803" severity error;
    assert SOL = '0' report "Error in test case #178/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #179/2803" severity error;
    assert SOR = '0' report "Error in test case #179/2803" severity error;
    assert SOL = '0' report "Error in test case #179/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #180/2803" severity error;
    assert SOR = '0' report "Error in test case #180/2803" severity error;
    assert SOL = '0' report "Error in test case #180/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #181/2803" severity error;
    assert SOR = '0' report "Error in test case #181/2803" severity error;
    assert SOL = '0' report "Error in test case #181/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #182/2803" severity error;
    assert SOR = '0' report "Error in test case #182/2803" severity error;
    assert SOL = '0' report "Error in test case #182/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #183/2803" severity error;
    assert SOR = '0' report "Error in test case #183/2803" severity error;
    assert SOL = '0' report "Error in test case #183/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #184/2803" severity error;
    assert SOR = '0' report "Error in test case #184/2803" severity error;
    assert SOL = '0' report "Error in test case #184/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #185/2803" severity error;
    assert SOR = '0' report "Error in test case #185/2803" severity error;
    assert SOL = '0' report "Error in test case #185/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #186/2803" severity error;
    assert SOR = '0' report "Error in test case #186/2803" severity error;
    assert SOL = '0' report "Error in test case #186/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #187/2803" severity error;
    assert SOR = '0' report "Error in test case #187/2803" severity error;
    assert SOL = '0' report "Error in test case #187/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #188/2803" severity error;
    assert SOR = '0' report "Error in test case #188/2803" severity error;
    assert SOL = '0' report "Error in test case #188/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #189/2803" severity error;
    assert SOR = '0' report "Error in test case #189/2803" severity error;
    assert SOL = '0' report "Error in test case #189/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #190/2803" severity error;
    assert SOR = '0' report "Error in test case #190/2803" severity error;
    assert SOL = '0' report "Error in test case #190/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #191/2803" severity error;
    assert SOR = '0' report "Error in test case #191/2803" severity error;
    assert SOL = '0' report "Error in test case #191/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #192/2803" severity error;
    assert SOR = '0' report "Error in test case #192/2803" severity error;
    assert SOL = '0' report "Error in test case #192/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #193/2803" severity error;
    assert SOR = '0' report "Error in test case #193/2803" severity error;
    assert SOL = '0' report "Error in test case #193/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #194/2803" severity error;
    assert SOR = '0' report "Error in test case #194/2803" severity error;
    assert SOL = '0' report "Error in test case #194/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #195/2803" severity error;
    assert SOR = '0' report "Error in test case #195/2803" severity error;
    assert SOL = '0' report "Error in test case #195/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #196/2803" severity error;
    assert SOR = '0' report "Error in test case #196/2803" severity error;
    assert SOL = '0' report "Error in test case #196/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #197/2803" severity error;
    assert SOR = '0' report "Error in test case #197/2803" severity error;
    assert SOL = '0' report "Error in test case #197/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #198/2803" severity error;
    assert SOR = '0' report "Error in test case #198/2803" severity error;
    assert SOL = '0' report "Error in test case #198/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #199/2803" severity error;
    assert SOR = '0' report "Error in test case #199/2803" severity error;
    assert SOL = '0' report "Error in test case #199/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #200/2803" severity error;
    assert SOR = '0' report "Error in test case #200/2803" severity error;
    assert SOL = '0' report "Error in test case #200/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #201/2803" severity error;
    assert SOR = '0' report "Error in test case #201/2803" severity error;
    assert SOL = '0' report "Error in test case #201/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #202/2803" severity error;
    assert SOR = '0' report "Error in test case #202/2803" severity error;
    assert SOL = '0' report "Error in test case #202/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #203/2803" severity error;
    assert SOR = '0' report "Error in test case #203/2803" severity error;
    assert SOL = '0' report "Error in test case #203/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #204/2803" severity error;
    assert SOR = '0' report "Error in test case #204/2803" severity error;
    assert SOL = '0' report "Error in test case #204/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #205/2803" severity error;
    assert SOR = '0' report "Error in test case #205/2803" severity error;
    assert SOL = '0' report "Error in test case #205/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #206/2803" severity error;
    assert SOR = '0' report "Error in test case #206/2803" severity error;
    assert SOL = '0' report "Error in test case #206/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #207/2803" severity error;
    assert SOR = '0' report "Error in test case #207/2803" severity error;
    assert SOL = '0' report "Error in test case #207/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #208/2803" severity error;
    assert SOR = '0' report "Error in test case #208/2803" severity error;
    assert SOL = '0' report "Error in test case #208/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #209/2803" severity error;
    assert SOR = '0' report "Error in test case #209/2803" severity error;
    assert SOL = '0' report "Error in test case #209/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #210/2803" severity error;
    assert SOR = '0' report "Error in test case #210/2803" severity error;
    assert SOL = '0' report "Error in test case #210/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #211/2803" severity error;
    assert SOR = '0' report "Error in test case #211/2803" severity error;
    assert SOL = '0' report "Error in test case #211/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #212/2803" severity error;
    assert SOR = '0' report "Error in test case #212/2803" severity error;
    assert SOL = '0' report "Error in test case #212/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #213/2803" severity error;
    assert SOR = '0' report "Error in test case #213/2803" severity error;
    assert SOL = '0' report "Error in test case #213/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #214/2803" severity error;
    assert SOR = '0' report "Error in test case #214/2803" severity error;
    assert SOL = '0' report "Error in test case #214/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #215/2803" severity error;
    assert SOR = '0' report "Error in test case #215/2803" severity error;
    assert SOL = '0' report "Error in test case #215/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #216/2803" severity error;
    assert SOR = '0' report "Error in test case #216/2803" severity error;
    assert SOL = '0' report "Error in test case #216/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #217/2803" severity error;
    assert SOR = '0' report "Error in test case #217/2803" severity error;
    assert SOL = '0' report "Error in test case #217/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #218/2803" severity error;
    assert SOR = '0' report "Error in test case #218/2803" severity error;
    assert SOL = '0' report "Error in test case #218/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #219/2803" severity error;
    assert SOR = '0' report "Error in test case #219/2803" severity error;
    assert SOL = '0' report "Error in test case #219/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #220/2803" severity error;
    assert SOR = '0' report "Error in test case #220/2803" severity error;
    assert SOL = '0' report "Error in test case #220/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #221/2803" severity error;
    assert SOR = '0' report "Error in test case #221/2803" severity error;
    assert SOL = '0' report "Error in test case #221/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #222/2803" severity error;
    assert SOR = '0' report "Error in test case #222/2803" severity error;
    assert SOL = '0' report "Error in test case #222/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #223/2803" severity error;
    assert SOR = '0' report "Error in test case #223/2803" severity error;
    assert SOL = '0' report "Error in test case #223/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #224/2803" severity error;
    assert SOR = '0' report "Error in test case #224/2803" severity error;
    assert SOL = '0' report "Error in test case #224/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #225/2803" severity error;
    assert SOR = '0' report "Error in test case #225/2803" severity error;
    assert SOL = '0' report "Error in test case #225/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #226/2803" severity error;
    assert SOR = '0' report "Error in test case #226/2803" severity error;
    assert SOL = '0' report "Error in test case #226/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #227/2803" severity error;
    assert SOR = '0' report "Error in test case #227/2803" severity error;
    assert SOL = '0' report "Error in test case #227/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #228/2803" severity error;
    assert SOR = '0' report "Error in test case #228/2803" severity error;
    assert SOL = '0' report "Error in test case #228/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #229/2803" severity error;
    assert SOR = '0' report "Error in test case #229/2803" severity error;
    assert SOL = '0' report "Error in test case #229/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #230/2803" severity error;
    assert SOR = '0' report "Error in test case #230/2803" severity error;
    assert SOL = '0' report "Error in test case #230/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #231/2803" severity error;
    assert SOR = '0' report "Error in test case #231/2803" severity error;
    assert SOL = '0' report "Error in test case #231/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #232/2803" severity error;
    assert SOR = '0' report "Error in test case #232/2803" severity error;
    assert SOL = '0' report "Error in test case #232/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #233/2803" severity error;
    assert SOR = '0' report "Error in test case #233/2803" severity error;
    assert SOL = '0' report "Error in test case #233/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #234/2803" severity error;
    assert SOR = '0' report "Error in test case #234/2803" severity error;
    assert SOL = '0' report "Error in test case #234/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #235/2803" severity error;
    assert SOR = '0' report "Error in test case #235/2803" severity error;
    assert SOL = '0' report "Error in test case #235/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #236/2803" severity error;
    assert SOR = '0' report "Error in test case #236/2803" severity error;
    assert SOL = '0' report "Error in test case #236/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #237/2803" severity error;
    assert SOR = '0' report "Error in test case #237/2803" severity error;
    assert SOL = '0' report "Error in test case #237/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #238/2803" severity error;
    assert SOR = '0' report "Error in test case #238/2803" severity error;
    assert SOL = '0' report "Error in test case #238/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #239/2803" severity error;
    assert SOR = '0' report "Error in test case #239/2803" severity error;
    assert SOL = '0' report "Error in test case #239/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #240/2803" severity error;
    assert SOR = '0' report "Error in test case #240/2803" severity error;
    assert SOL = '0' report "Error in test case #240/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #241/2803" severity error;
    assert SOR = '0' report "Error in test case #241/2803" severity error;
    assert SOL = '0' report "Error in test case #241/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #242/2803" severity error;
    assert SOR = '0' report "Error in test case #242/2803" severity error;
    assert SOL = '0' report "Error in test case #242/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #243/2803" severity error;
    assert SOR = '0' report "Error in test case #243/2803" severity error;
    assert SOL = '0' report "Error in test case #243/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #244/2803" severity error;
    assert SOR = '0' report "Error in test case #244/2803" severity error;
    assert SOL = '0' report "Error in test case #244/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #245/2803" severity error;
    assert SOR = '0' report "Error in test case #245/2803" severity error;
    assert SOL = '0' report "Error in test case #245/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #246/2803" severity error;
    assert SOR = '0' report "Error in test case #246/2803" severity error;
    assert SOL = '0' report "Error in test case #246/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #247/2803" severity error;
    assert SOR = '0' report "Error in test case #247/2803" severity error;
    assert SOL = '0' report "Error in test case #247/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #248/2803" severity error;
    assert SOR = '0' report "Error in test case #248/2803" severity error;
    assert SOL = '0' report "Error in test case #248/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #249/2803" severity error;
    assert SOR = '0' report "Error in test case #249/2803" severity error;
    assert SOL = '0' report "Error in test case #249/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #250/2803" severity error;
    assert SOR = '0' report "Error in test case #250/2803" severity error;
    assert SOL = '0' report "Error in test case #250/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #251/2803" severity error;
    assert SOR = '0' report "Error in test case #251/2803" severity error;
    assert SOL = '0' report "Error in test case #251/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #252/2803" severity error;
    assert SOR = '0' report "Error in test case #252/2803" severity error;
    assert SOL = '0' report "Error in test case #252/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #253/2803" severity error;
    assert SOR = '0' report "Error in test case #253/2803" severity error;
    assert SOL = '0' report "Error in test case #253/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #254/2803" severity error;
    assert SOR = '0' report "Error in test case #254/2803" severity error;
    assert SOL = '0' report "Error in test case #254/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #255/2803" severity error;
    assert SOR = '0' report "Error in test case #255/2803" severity error;
    assert SOL = '0' report "Error in test case #255/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #256/2803" severity error;
    assert SOR = '0' report "Error in test case #256/2803" severity error;
    assert SOL = '0' report "Error in test case #256/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #257/2803" severity error;
    assert SOR = '0' report "Error in test case #257/2803" severity error;
    assert SOL = '0' report "Error in test case #257/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #258/2803" severity error;
    assert SOR = '0' report "Error in test case #258/2803" severity error;
    assert SOL = '0' report "Error in test case #258/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #259/2803" severity error;
    assert SOR = '0' report "Error in test case #259/2803" severity error;
    assert SOL = '0' report "Error in test case #259/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #260/2803" severity error;
    assert SOR = '0' report "Error in test case #260/2803" severity error;
    assert SOL = '0' report "Error in test case #260/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #261/2803" severity error;
    assert SOR = '0' report "Error in test case #261/2803" severity error;
    assert SOL = '0' report "Error in test case #261/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #262/2803" severity error;
    assert SOR = '0' report "Error in test case #262/2803" severity error;
    assert SOL = '0' report "Error in test case #262/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #263/2803" severity error;
    assert SOR = '0' report "Error in test case #263/2803" severity error;
    assert SOL = '0' report "Error in test case #263/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #264/2803" severity error;
    assert SOR = '0' report "Error in test case #264/2803" severity error;
    assert SOL = '0' report "Error in test case #264/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #265/2803" severity error;
    assert SOR = '0' report "Error in test case #265/2803" severity error;
    assert SOL = '0' report "Error in test case #265/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #266/2803" severity error;
    assert SOR = '0' report "Error in test case #266/2803" severity error;
    assert SOL = '0' report "Error in test case #266/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #267/2803" severity error;
    assert SOR = '0' report "Error in test case #267/2803" severity error;
    assert SOL = '0' report "Error in test case #267/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #268/2803" severity error;
    assert SOR = '0' report "Error in test case #268/2803" severity error;
    assert SOL = '0' report "Error in test case #268/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #269/2803" severity error;
    assert SOR = '0' report "Error in test case #269/2803" severity error;
    assert SOL = '0' report "Error in test case #269/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #270/2803" severity error;
    assert SOR = '0' report "Error in test case #270/2803" severity error;
    assert SOL = '0' report "Error in test case #270/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #271/2803" severity error;
    assert SOR = '0' report "Error in test case #271/2803" severity error;
    assert SOL = '0' report "Error in test case #271/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #272/2803" severity error;
    assert SOR = '1' report "Error in test case #272/2803" severity error;
    assert SOL = '1' report "Error in test case #272/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #273/2803" severity error;
    assert SOR = '1' report "Error in test case #273/2803" severity error;
    assert SOL = '1' report "Error in test case #273/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #274/2803" severity error;
    assert SOR = '1' report "Error in test case #274/2803" severity error;
    assert SOL = '1' report "Error in test case #274/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #275/2803" severity error;
    assert SOR = '1' report "Error in test case #275/2803" severity error;
    assert SOL = '1' report "Error in test case #275/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #276/2803" severity error;
    assert SOR = '1' report "Error in test case #276/2803" severity error;
    assert SOL = '1' report "Error in test case #276/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #277/2803" severity error;
    assert SOR = '1' report "Error in test case #277/2803" severity error;
    assert SOL = '1' report "Error in test case #277/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #278/2803" severity error;
    assert SOR = '1' report "Error in test case #278/2803" severity error;
    assert SOL = '1' report "Error in test case #278/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #279/2803" severity error;
    assert SOR = '1' report "Error in test case #279/2803" severity error;
    assert SOL = '1' report "Error in test case #279/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #280/2803" severity error;
    assert SOR = '1' report "Error in test case #280/2803" severity error;
    assert SOL = '1' report "Error in test case #280/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #281/2803" severity error;
    assert SOR = '1' report "Error in test case #281/2803" severity error;
    assert SOL = '1' report "Error in test case #281/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #282/2803" severity error;
    assert SOR = '1' report "Error in test case #282/2803" severity error;
    assert SOL = '1' report "Error in test case #282/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #283/2803" severity error;
    assert SOR = '1' report "Error in test case #283/2803" severity error;
    assert SOL = '1' report "Error in test case #283/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #284/2803" severity error;
    assert SOR = '1' report "Error in test case #284/2803" severity error;
    assert SOL = '1' report "Error in test case #284/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #285/2803" severity error;
    assert SOR = '1' report "Error in test case #285/2803" severity error;
    assert SOL = '1' report "Error in test case #285/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #286/2803" severity error;
    assert SOR = '1' report "Error in test case #286/2803" severity error;
    assert SOL = '1' report "Error in test case #286/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #287/2803" severity error;
    assert SOR = '1' report "Error in test case #287/2803" severity error;
    assert SOL = '1' report "Error in test case #287/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #288/2803" severity error;
    assert SOR = '1' report "Error in test case #288/2803" severity error;
    assert SOL = '1' report "Error in test case #288/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #289/2803" severity error;
    assert SOR = '1' report "Error in test case #289/2803" severity error;
    assert SOL = '1' report "Error in test case #289/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #290/2803" severity error;
    assert SOR = '1' report "Error in test case #290/2803" severity error;
    assert SOL = '1' report "Error in test case #290/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #291/2803" severity error;
    assert SOR = '1' report "Error in test case #291/2803" severity error;
    assert SOL = '1' report "Error in test case #291/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #292/2803" severity error;
    assert SOR = '1' report "Error in test case #292/2803" severity error;
    assert SOL = '1' report "Error in test case #292/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #293/2803" severity error;
    assert SOR = '1' report "Error in test case #293/2803" severity error;
    assert SOL = '1' report "Error in test case #293/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #294/2803" severity error;
    assert SOR = '1' report "Error in test case #294/2803" severity error;
    assert SOL = '1' report "Error in test case #294/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #295/2803" severity error;
    assert SOR = '1' report "Error in test case #295/2803" severity error;
    assert SOL = '1' report "Error in test case #295/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #296/2803" severity error;
    assert SOR = '1' report "Error in test case #296/2803" severity error;
    assert SOL = '1' report "Error in test case #296/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #297/2803" severity error;
    assert SOR = '1' report "Error in test case #297/2803" severity error;
    assert SOL = '1' report "Error in test case #297/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #298/2803" severity error;
    assert SOR = '1' report "Error in test case #298/2803" severity error;
    assert SOL = '1' report "Error in test case #298/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #299/2803" severity error;
    assert SOR = '1' report "Error in test case #299/2803" severity error;
    assert SOL = '1' report "Error in test case #299/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #300/2803" severity error;
    assert SOR = '1' report "Error in test case #300/2803" severity error;
    assert SOL = '1' report "Error in test case #300/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #301/2803" severity error;
    assert SOR = '1' report "Error in test case #301/2803" severity error;
    assert SOL = '1' report "Error in test case #301/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #302/2803" severity error;
    assert SOR = '1' report "Error in test case #302/2803" severity error;
    assert SOL = '1' report "Error in test case #302/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #303/2803" severity error;
    assert SOR = '1' report "Error in test case #303/2803" severity error;
    assert SOL = '1' report "Error in test case #303/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #304/2803" severity error;
    assert SOR = '1' report "Error in test case #304/2803" severity error;
    assert SOL = '1' report "Error in test case #304/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #305/2803" severity error;
    assert SOR = '1' report "Error in test case #305/2803" severity error;
    assert SOL = '1' report "Error in test case #305/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #306/2803" severity error;
    assert SOR = '1' report "Error in test case #306/2803" severity error;
    assert SOL = '1' report "Error in test case #306/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #307/2803" severity error;
    assert SOR = '1' report "Error in test case #307/2803" severity error;
    assert SOL = '1' report "Error in test case #307/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #308/2803" severity error;
    assert SOR = '1' report "Error in test case #308/2803" severity error;
    assert SOL = '1' report "Error in test case #308/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #309/2803" severity error;
    assert SOR = '1' report "Error in test case #309/2803" severity error;
    assert SOL = '1' report "Error in test case #309/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #310/2803" severity error;
    assert SOR = '1' report "Error in test case #310/2803" severity error;
    assert SOL = '1' report "Error in test case #310/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #311/2803" severity error;
    assert SOR = '1' report "Error in test case #311/2803" severity error;
    assert SOL = '1' report "Error in test case #311/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #312/2803" severity error;
    assert SOR = '1' report "Error in test case #312/2803" severity error;
    assert SOL = '1' report "Error in test case #312/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #313/2803" severity error;
    assert SOR = '1' report "Error in test case #313/2803" severity error;
    assert SOL = '1' report "Error in test case #313/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #314/2803" severity error;
    assert SOR = '1' report "Error in test case #314/2803" severity error;
    assert SOL = '1' report "Error in test case #314/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #315/2803" severity error;
    assert SOR = '1' report "Error in test case #315/2803" severity error;
    assert SOL = '1' report "Error in test case #315/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #316/2803" severity error;
    assert SOR = '1' report "Error in test case #316/2803" severity error;
    assert SOL = '1' report "Error in test case #316/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #317/2803" severity error;
    assert SOR = '1' report "Error in test case #317/2803" severity error;
    assert SOL = '1' report "Error in test case #317/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #318/2803" severity error;
    assert SOR = '1' report "Error in test case #318/2803" severity error;
    assert SOL = '1' report "Error in test case #318/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #319/2803" severity error;
    assert SOR = '1' report "Error in test case #319/2803" severity error;
    assert SOL = '1' report "Error in test case #319/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #320/2803" severity error;
    assert SOR = '1' report "Error in test case #320/2803" severity error;
    assert SOL = '1' report "Error in test case #320/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #321/2803" severity error;
    assert SOR = '1' report "Error in test case #321/2803" severity error;
    assert SOL = '1' report "Error in test case #321/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #322/2803" severity error;
    assert SOR = '1' report "Error in test case #322/2803" severity error;
    assert SOL = '1' report "Error in test case #322/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #323/2803" severity error;
    assert SOR = '1' report "Error in test case #323/2803" severity error;
    assert SOL = '1' report "Error in test case #323/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #324/2803" severity error;
    assert SOR = '1' report "Error in test case #324/2803" severity error;
    assert SOL = '1' report "Error in test case #324/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #325/2803" severity error;
    assert SOR = '1' report "Error in test case #325/2803" severity error;
    assert SOL = '1' report "Error in test case #325/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #326/2803" severity error;
    assert SOR = '1' report "Error in test case #326/2803" severity error;
    assert SOL = '1' report "Error in test case #326/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #327/2803" severity error;
    assert SOR = '1' report "Error in test case #327/2803" severity error;
    assert SOL = '1' report "Error in test case #327/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #328/2803" severity error;
    assert SOR = '1' report "Error in test case #328/2803" severity error;
    assert SOL = '1' report "Error in test case #328/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #329/2803" severity error;
    assert SOR = '1' report "Error in test case #329/2803" severity error;
    assert SOL = '1' report "Error in test case #329/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #330/2803" severity error;
    assert SOR = '1' report "Error in test case #330/2803" severity error;
    assert SOL = '1' report "Error in test case #330/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #331/2803" severity error;
    assert SOR = '1' report "Error in test case #331/2803" severity error;
    assert SOL = '1' report "Error in test case #331/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #332/2803" severity error;
    assert SOR = '1' report "Error in test case #332/2803" severity error;
    assert SOL = '1' report "Error in test case #332/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #333/2803" severity error;
    assert SOR = '1' report "Error in test case #333/2803" severity error;
    assert SOL = '1' report "Error in test case #333/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #334/2803" severity error;
    assert SOR = '1' report "Error in test case #334/2803" severity error;
    assert SOL = '1' report "Error in test case #334/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #335/2803" severity error;
    assert SOR = '1' report "Error in test case #335/2803" severity error;
    assert SOL = '1' report "Error in test case #335/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #336/2803" severity error;
    assert SOR = '1' report "Error in test case #336/2803" severity error;
    assert SOL = '1' report "Error in test case #336/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #337/2803" severity error;
    assert SOR = '1' report "Error in test case #337/2803" severity error;
    assert SOL = '1' report "Error in test case #337/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #338/2803" severity error;
    assert SOR = '1' report "Error in test case #338/2803" severity error;
    assert SOL = '1' report "Error in test case #338/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #339/2803" severity error;
    assert SOR = '1' report "Error in test case #339/2803" severity error;
    assert SOL = '1' report "Error in test case #339/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #340/2803" severity error;
    assert SOR = '1' report "Error in test case #340/2803" severity error;
    assert SOL = '1' report "Error in test case #340/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #341/2803" severity error;
    assert SOR = '1' report "Error in test case #341/2803" severity error;
    assert SOL = '1' report "Error in test case #341/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #342/2803" severity error;
    assert SOR = '1' report "Error in test case #342/2803" severity error;
    assert SOL = '1' report "Error in test case #342/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #343/2803" severity error;
    assert SOR = '1' report "Error in test case #343/2803" severity error;
    assert SOL = '1' report "Error in test case #343/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #344/2803" severity error;
    assert SOR = '1' report "Error in test case #344/2803" severity error;
    assert SOL = '1' report "Error in test case #344/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #345/2803" severity error;
    assert SOR = '1' report "Error in test case #345/2803" severity error;
    assert SOL = '1' report "Error in test case #345/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #346/2803" severity error;
    assert SOR = '1' report "Error in test case #346/2803" severity error;
    assert SOL = '1' report "Error in test case #346/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #347/2803" severity error;
    assert SOR = '1' report "Error in test case #347/2803" severity error;
    assert SOL = '1' report "Error in test case #347/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #348/2803" severity error;
    assert SOR = '1' report "Error in test case #348/2803" severity error;
    assert SOL = '1' report "Error in test case #348/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #349/2803" severity error;
    assert SOR = '1' report "Error in test case #349/2803" severity error;
    assert SOL = '1' report "Error in test case #349/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #350/2803" severity error;
    assert SOR = '1' report "Error in test case #350/2803" severity error;
    assert SOL = '1' report "Error in test case #350/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #351/2803" severity error;
    assert SOR = '1' report "Error in test case #351/2803" severity error;
    assert SOL = '1' report "Error in test case #351/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #352/2803" severity error;
    assert SOR = '1' report "Error in test case #352/2803" severity error;
    assert SOL = '1' report "Error in test case #352/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #353/2803" severity error;
    assert SOR = '1' report "Error in test case #353/2803" severity error;
    assert SOL = '1' report "Error in test case #353/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #354/2803" severity error;
    assert SOR = '1' report "Error in test case #354/2803" severity error;
    assert SOL = '1' report "Error in test case #354/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #355/2803" severity error;
    assert SOR = '1' report "Error in test case #355/2803" severity error;
    assert SOL = '1' report "Error in test case #355/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #356/2803" severity error;
    assert SOR = '1' report "Error in test case #356/2803" severity error;
    assert SOL = '1' report "Error in test case #356/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #357/2803" severity error;
    assert SOR = '1' report "Error in test case #357/2803" severity error;
    assert SOL = '1' report "Error in test case #357/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #358/2803" severity error;
    assert SOR = '1' report "Error in test case #358/2803" severity error;
    assert SOL = '1' report "Error in test case #358/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #359/2803" severity error;
    assert SOR = '1' report "Error in test case #359/2803" severity error;
    assert SOL = '1' report "Error in test case #359/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #360/2803" severity error;
    assert SOR = '1' report "Error in test case #360/2803" severity error;
    assert SOL = '1' report "Error in test case #360/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #361/2803" severity error;
    assert SOR = '1' report "Error in test case #361/2803" severity error;
    assert SOL = '1' report "Error in test case #361/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #362/2803" severity error;
    assert SOR = '1' report "Error in test case #362/2803" severity error;
    assert SOL = '1' report "Error in test case #362/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #363/2803" severity error;
    assert SOR = '1' report "Error in test case #363/2803" severity error;
    assert SOL = '1' report "Error in test case #363/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #364/2803" severity error;
    assert SOR = '1' report "Error in test case #364/2803" severity error;
    assert SOL = '1' report "Error in test case #364/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #365/2803" severity error;
    assert SOR = '1' report "Error in test case #365/2803" severity error;
    assert SOL = '1' report "Error in test case #365/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #366/2803" severity error;
    assert SOR = '1' report "Error in test case #366/2803" severity error;
    assert SOL = '1' report "Error in test case #366/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #367/2803" severity error;
    assert SOR = '1' report "Error in test case #367/2803" severity error;
    assert SOL = '1' report "Error in test case #367/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #368/2803" severity error;
    assert SOR = '1' report "Error in test case #368/2803" severity error;
    assert SOL = '1' report "Error in test case #368/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #369/2803" severity error;
    assert SOR = '1' report "Error in test case #369/2803" severity error;
    assert SOL = '1' report "Error in test case #369/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #370/2803" severity error;
    assert SOR = '1' report "Error in test case #370/2803" severity error;
    assert SOL = '1' report "Error in test case #370/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #371/2803" severity error;
    assert SOR = '1' report "Error in test case #371/2803" severity error;
    assert SOL = '1' report "Error in test case #371/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #372/2803" severity error;
    assert SOR = '1' report "Error in test case #372/2803" severity error;
    assert SOL = '1' report "Error in test case #372/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #373/2803" severity error;
    assert SOR = '1' report "Error in test case #373/2803" severity error;
    assert SOL = '1' report "Error in test case #373/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #374/2803" severity error;
    assert SOR = '1' report "Error in test case #374/2803" severity error;
    assert SOL = '1' report "Error in test case #374/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #375/2803" severity error;
    assert SOR = '1' report "Error in test case #375/2803" severity error;
    assert SOL = '1' report "Error in test case #375/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #376/2803" severity error;
    assert SOR = '1' report "Error in test case #376/2803" severity error;
    assert SOL = '1' report "Error in test case #376/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #377/2803" severity error;
    assert SOR = '1' report "Error in test case #377/2803" severity error;
    assert SOL = '1' report "Error in test case #377/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #378/2803" severity error;
    assert SOR = '1' report "Error in test case #378/2803" severity error;
    assert SOL = '1' report "Error in test case #378/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #379/2803" severity error;
    assert SOR = '1' report "Error in test case #379/2803" severity error;
    assert SOL = '1' report "Error in test case #379/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #380/2803" severity error;
    assert SOR = '1' report "Error in test case #380/2803" severity error;
    assert SOL = '1' report "Error in test case #380/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #381/2803" severity error;
    assert SOR = '1' report "Error in test case #381/2803" severity error;
    assert SOL = '1' report "Error in test case #381/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #382/2803" severity error;
    assert SOR = '1' report "Error in test case #382/2803" severity error;
    assert SOL = '1' report "Error in test case #382/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #383/2803" severity error;
    assert SOR = '0' report "Error in test case #383/2803" severity error;
    assert SOL = '0' report "Error in test case #383/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #384/2803" severity error;
    assert SOR = '0' report "Error in test case #384/2803" severity error;
    assert SOL = '0' report "Error in test case #384/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #385/2803" severity error;
    assert SOR = '0' report "Error in test case #385/2803" severity error;
    assert SOL = '0' report "Error in test case #385/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #386/2803" severity error;
    assert SOR = '0' report "Error in test case #386/2803" severity error;
    assert SOL = '0' report "Error in test case #386/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #387/2803" severity error;
    assert SOR = '0' report "Error in test case #387/2803" severity error;
    assert SOL = '0' report "Error in test case #387/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #388/2803" severity error;
    assert SOR = '0' report "Error in test case #388/2803" severity error;
    assert SOL = '0' report "Error in test case #388/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #389/2803" severity error;
    assert SOR = '0' report "Error in test case #389/2803" severity error;
    assert SOL = '0' report "Error in test case #389/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #390/2803" severity error;
    assert SOR = '0' report "Error in test case #390/2803" severity error;
    assert SOL = '0' report "Error in test case #390/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #391/2803" severity error;
    assert SOR = '0' report "Error in test case #391/2803" severity error;
    assert SOL = '0' report "Error in test case #391/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #392/2803" severity error;
    assert SOR = '0' report "Error in test case #392/2803" severity error;
    assert SOL = '0' report "Error in test case #392/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #393/2803" severity error;
    assert SOR = '0' report "Error in test case #393/2803" severity error;
    assert SOL = '0' report "Error in test case #393/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #394/2803" severity error;
    assert SOR = '0' report "Error in test case #394/2803" severity error;
    assert SOL = '0' report "Error in test case #394/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #395/2803" severity error;
    assert SOR = '0' report "Error in test case #395/2803" severity error;
    assert SOL = '0' report "Error in test case #395/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #396/2803" severity error;
    assert SOR = '0' report "Error in test case #396/2803" severity error;
    assert SOL = '0' report "Error in test case #396/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #397/2803" severity error;
    assert SOR = '0' report "Error in test case #397/2803" severity error;
    assert SOL = '0' report "Error in test case #397/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #398/2803" severity error;
    assert SOR = '0' report "Error in test case #398/2803" severity error;
    assert SOL = '0' report "Error in test case #398/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #399/2803" severity error;
    assert SOR = '0' report "Error in test case #399/2803" severity error;
    assert SOL = '0' report "Error in test case #399/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #400/2803" severity error;
    assert SOR = '0' report "Error in test case #400/2803" severity error;
    assert SOL = '0' report "Error in test case #400/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #401/2803" severity error;
    assert SOR = '0' report "Error in test case #401/2803" severity error;
    assert SOL = '0' report "Error in test case #401/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #402/2803" severity error;
    assert SOR = '0' report "Error in test case #402/2803" severity error;
    assert SOL = '0' report "Error in test case #402/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "000";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #403/2803" severity error;
    assert SOR = '0' report "Error in test case #403/2803" severity error;
    assert SOL = '0' report "Error in test case #403/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #404/2803" severity error;
    assert SOR = '0' report "Error in test case #404/2803" severity error;
    assert SOL = '0' report "Error in test case #404/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #405/2803" severity error;
    assert SOR = '0' report "Error in test case #405/2803" severity error;
    assert SOL = '0' report "Error in test case #405/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #406/2803" severity error;
    assert SOR = '0' report "Error in test case #406/2803" severity error;
    assert SOL = '0' report "Error in test case #406/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #407/2803" severity error;
    assert SOR = '0' report "Error in test case #407/2803" severity error;
    assert SOL = '0' report "Error in test case #407/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #408/2803" severity error;
    assert SOR = '0' report "Error in test case #408/2803" severity error;
    assert SOL = '1' report "Error in test case #408/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #409/2803" severity error;
    assert SOR = '0' report "Error in test case #409/2803" severity error;
    assert SOL = '1' report "Error in test case #409/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #410/2803" severity error;
    assert SOR = '0' report "Error in test case #410/2803" severity error;
    assert SOL = '1' report "Error in test case #410/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #411/2803" severity error;
    assert SOR = '0' report "Error in test case #411/2803" severity error;
    assert SOL = '1' report "Error in test case #411/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #412/2803" severity error;
    assert SOR = '0' report "Error in test case #412/2803" severity error;
    assert SOL = '1' report "Error in test case #412/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #413/2803" severity error;
    assert SOR = '0' report "Error in test case #413/2803" severity error;
    assert SOL = '1' report "Error in test case #413/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #414/2803" severity error;
    assert SOR = '0' report "Error in test case #414/2803" severity error;
    assert SOL = '1' report "Error in test case #414/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #415/2803" severity error;
    assert SOR = '0' report "Error in test case #415/2803" severity error;
    assert SOL = '1' report "Error in test case #415/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #416/2803" severity error;
    assert SOR = '0' report "Error in test case #416/2803" severity error;
    assert SOL = '0' report "Error in test case #416/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #417/2803" severity error;
    assert SOR = '0' report "Error in test case #417/2803" severity error;
    assert SOL = '0' report "Error in test case #417/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #418/2803" severity error;
    assert SOR = '0' report "Error in test case #418/2803" severity error;
    assert SOL = '0' report "Error in test case #418/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #419/2803" severity error;
    assert SOR = '0' report "Error in test case #419/2803" severity error;
    assert SOL = '0' report "Error in test case #419/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #420/2803" severity error;
    assert SOR = '0' report "Error in test case #420/2803" severity error;
    assert SOL = '0' report "Error in test case #420/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #421/2803" severity error;
    assert SOR = '0' report "Error in test case #421/2803" severity error;
    assert SOL = '0' report "Error in test case #421/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #422/2803" severity error;
    assert SOR = '0' report "Error in test case #422/2803" severity error;
    assert SOL = '0' report "Error in test case #422/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #423/2803" severity error;
    assert SOR = '0' report "Error in test case #423/2803" severity error;
    assert SOL = '0' report "Error in test case #423/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00100000" report "Error in test case #424/2803" severity error;
    assert SOR = '0' report "Error in test case #424/2803" severity error;
    assert SOL = '0' report "Error in test case #424/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00100000" report "Error in test case #425/2803" severity error;
    assert SOR = '0' report "Error in test case #425/2803" severity error;
    assert SOL = '0' report "Error in test case #425/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00100000" report "Error in test case #426/2803" severity error;
    assert SOR = '0' report "Error in test case #426/2803" severity error;
    assert SOL = '0' report "Error in test case #426/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00100000" report "Error in test case #427/2803" severity error;
    assert SOR = '0' report "Error in test case #427/2803" severity error;
    assert SOL = '0' report "Error in test case #427/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00100000" report "Error in test case #428/2803" severity error;
    assert SOR = '0' report "Error in test case #428/2803" severity error;
    assert SOL = '0' report "Error in test case #428/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00100000" report "Error in test case #429/2803" severity error;
    assert SOR = '0' report "Error in test case #429/2803" severity error;
    assert SOL = '0' report "Error in test case #429/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00100000" report "Error in test case #430/2803" severity error;
    assert SOR = '0' report "Error in test case #430/2803" severity error;
    assert SOL = '0' report "Error in test case #430/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00100000" report "Error in test case #431/2803" severity error;
    assert SOR = '0' report "Error in test case #431/2803" severity error;
    assert SOL = '0' report "Error in test case #431/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010000" report "Error in test case #432/2803" severity error;
    assert SOR = '0' report "Error in test case #432/2803" severity error;
    assert SOL = '1' report "Error in test case #432/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010000" report "Error in test case #433/2803" severity error;
    assert SOR = '0' report "Error in test case #433/2803" severity error;
    assert SOL = '1' report "Error in test case #433/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010000" report "Error in test case #434/2803" severity error;
    assert SOR = '0' report "Error in test case #434/2803" severity error;
    assert SOL = '1' report "Error in test case #434/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010000" report "Error in test case #435/2803" severity error;
    assert SOR = '0' report "Error in test case #435/2803" severity error;
    assert SOL = '1' report "Error in test case #435/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010000" report "Error in test case #436/2803" severity error;
    assert SOR = '0' report "Error in test case #436/2803" severity error;
    assert SOL = '1' report "Error in test case #436/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010000" report "Error in test case #437/2803" severity error;
    assert SOR = '0' report "Error in test case #437/2803" severity error;
    assert SOL = '1' report "Error in test case #437/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010000" report "Error in test case #438/2803" severity error;
    assert SOR = '0' report "Error in test case #438/2803" severity error;
    assert SOL = '1' report "Error in test case #438/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010000" report "Error in test case #439/2803" severity error;
    assert SOR = '0' report "Error in test case #439/2803" severity error;
    assert SOL = '1' report "Error in test case #439/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01001000" report "Error in test case #440/2803" severity error;
    assert SOR = '0' report "Error in test case #440/2803" severity error;
    assert SOL = '0' report "Error in test case #440/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01001000" report "Error in test case #441/2803" severity error;
    assert SOR = '0' report "Error in test case #441/2803" severity error;
    assert SOL = '0' report "Error in test case #441/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01001000" report "Error in test case #442/2803" severity error;
    assert SOR = '0' report "Error in test case #442/2803" severity error;
    assert SOL = '0' report "Error in test case #442/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #443/2803" severity error;
    assert SOR = '0' report "Error in test case #443/2803" severity error;
    assert SOL = '0' report "Error in test case #443/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #444/2803" severity error;
    assert SOR = '0' report "Error in test case #444/2803" severity error;
    assert SOL = '0' report "Error in test case #444/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #445/2803" severity error;
    assert SOR = '0' report "Error in test case #445/2803" severity error;
    assert SOL = '0' report "Error in test case #445/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #446/2803" severity error;
    assert SOR = '0' report "Error in test case #446/2803" severity error;
    assert SOL = '0' report "Error in test case #446/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #447/2803" severity error;
    assert SOR = '0' report "Error in test case #447/2803" severity error;
    assert SOL = '0' report "Error in test case #447/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #448/2803" severity error;
    assert SOR = '0' report "Error in test case #448/2803" severity error;
    assert SOL = '1' report "Error in test case #448/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #449/2803" severity error;
    assert SOR = '0' report "Error in test case #449/2803" severity error;
    assert SOL = '1' report "Error in test case #449/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #450/2803" severity error;
    assert SOR = '0' report "Error in test case #450/2803" severity error;
    assert SOL = '1' report "Error in test case #450/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #451/2803" severity error;
    assert SOR = '0' report "Error in test case #451/2803" severity error;
    assert SOL = '1' report "Error in test case #451/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #452/2803" severity error;
    assert SOR = '0' report "Error in test case #452/2803" severity error;
    assert SOL = '1' report "Error in test case #452/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #453/2803" severity error;
    assert SOR = '0' report "Error in test case #453/2803" severity error;
    assert SOL = '1' report "Error in test case #453/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #454/2803" severity error;
    assert SOR = '0' report "Error in test case #454/2803" severity error;
    assert SOL = '1' report "Error in test case #454/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #455/2803" severity error;
    assert SOR = '0' report "Error in test case #455/2803" severity error;
    assert SOL = '1' report "Error in test case #455/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #456/2803" severity error;
    assert SOR = '0' report "Error in test case #456/2803" severity error;
    assert SOL = '0' report "Error in test case #456/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #457/2803" severity error;
    assert SOR = '0' report "Error in test case #457/2803" severity error;
    assert SOL = '0' report "Error in test case #457/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #458/2803" severity error;
    assert SOR = '0' report "Error in test case #458/2803" severity error;
    assert SOL = '0' report "Error in test case #458/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #459/2803" severity error;
    assert SOR = '0' report "Error in test case #459/2803" severity error;
    assert SOL = '0' report "Error in test case #459/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #460/2803" severity error;
    assert SOR = '0' report "Error in test case #460/2803" severity error;
    assert SOL = '0' report "Error in test case #460/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #461/2803" severity error;
    assert SOR = '0' report "Error in test case #461/2803" severity error;
    assert SOL = '0' report "Error in test case #461/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #462/2803" severity error;
    assert SOR = '0' report "Error in test case #462/2803" severity error;
    assert SOL = '0' report "Error in test case #462/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01000000" report "Error in test case #463/2803" severity error;
    assert SOR = '0' report "Error in test case #463/2803" severity error;
    assert SOL = '0' report "Error in test case #463/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10100000" report "Error in test case #464/2803" severity error;
    assert SOR = '0' report "Error in test case #464/2803" severity error;
    assert SOL = '1' report "Error in test case #464/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10100000" report "Error in test case #465/2803" severity error;
    assert SOR = '0' report "Error in test case #465/2803" severity error;
    assert SOL = '1' report "Error in test case #465/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10100000" report "Error in test case #466/2803" severity error;
    assert SOR = '0' report "Error in test case #466/2803" severity error;
    assert SOL = '1' report "Error in test case #466/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10100000" report "Error in test case #467/2803" severity error;
    assert SOR = '0' report "Error in test case #467/2803" severity error;
    assert SOL = '1' report "Error in test case #467/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10100000" report "Error in test case #468/2803" severity error;
    assert SOR = '0' report "Error in test case #468/2803" severity error;
    assert SOL = '1' report "Error in test case #468/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10100000" report "Error in test case #469/2803" severity error;
    assert SOR = '0' report "Error in test case #469/2803" severity error;
    assert SOL = '1' report "Error in test case #469/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10100000" report "Error in test case #470/2803" severity error;
    assert SOR = '0' report "Error in test case #470/2803" severity error;
    assert SOL = '1' report "Error in test case #470/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10100000" report "Error in test case #471/2803" severity error;
    assert SOR = '0' report "Error in test case #471/2803" severity error;
    assert SOL = '1' report "Error in test case #471/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #472/2803" severity error;
    assert SOR = '1' report "Error in test case #472/2803" severity error;
    assert SOL = '1' report "Error in test case #472/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #473/2803" severity error;
    assert SOR = '1' report "Error in test case #473/2803" severity error;
    assert SOL = '1' report "Error in test case #473/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #474/2803" severity error;
    assert SOR = '1' report "Error in test case #474/2803" severity error;
    assert SOL = '1' report "Error in test case #474/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #475/2803" severity error;
    assert SOR = '1' report "Error in test case #475/2803" severity error;
    assert SOL = '1' report "Error in test case #475/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #476/2803" severity error;
    assert SOR = '1' report "Error in test case #476/2803" severity error;
    assert SOL = '1' report "Error in test case #476/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #477/2803" severity error;
    assert SOR = '1' report "Error in test case #477/2803" severity error;
    assert SOL = '1' report "Error in test case #477/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #478/2803" severity error;
    assert SOR = '1' report "Error in test case #478/2803" severity error;
    assert SOL = '1' report "Error in test case #478/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #479/2803" severity error;
    assert SOR = '1' report "Error in test case #479/2803" severity error;
    assert SOL = '1' report "Error in test case #479/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #480/2803" severity error;
    assert SOR = '1' report "Error in test case #480/2803" severity error;
    assert SOL = '0' report "Error in test case #480/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #481/2803" severity error;
    assert SOR = '1' report "Error in test case #481/2803" severity error;
    assert SOL = '0' report "Error in test case #481/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #482/2803" severity error;
    assert SOR = '1' report "Error in test case #482/2803" severity error;
    assert SOL = '0' report "Error in test case #482/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #483/2803" severity error;
    assert SOR = '1' report "Error in test case #483/2803" severity error;
    assert SOL = '0' report "Error in test case #483/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #484/2803" severity error;
    assert SOR = '1' report "Error in test case #484/2803" severity error;
    assert SOL = '0' report "Error in test case #484/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #485/2803" severity error;
    assert SOR = '1' report "Error in test case #485/2803" severity error;
    assert SOL = '0' report "Error in test case #485/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #486/2803" severity error;
    assert SOR = '1' report "Error in test case #486/2803" severity error;
    assert SOL = '0' report "Error in test case #486/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #487/2803" severity error;
    assert SOR = '1' report "Error in test case #487/2803" severity error;
    assert SOL = '0' report "Error in test case #487/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #488/2803" severity error;
    assert SOR = '1' report "Error in test case #488/2803" severity error;
    assert SOL = '0' report "Error in test case #488/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #489/2803" severity error;
    assert SOR = '1' report "Error in test case #489/2803" severity error;
    assert SOL = '0' report "Error in test case #489/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #490/2803" severity error;
    assert SOR = '1' report "Error in test case #490/2803" severity error;
    assert SOL = '0' report "Error in test case #490/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #491/2803" severity error;
    assert SOR = '1' report "Error in test case #491/2803" severity error;
    assert SOL = '0' report "Error in test case #491/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #492/2803" severity error;
    assert SOR = '1' report "Error in test case #492/2803" severity error;
    assert SOL = '0' report "Error in test case #492/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #493/2803" severity error;
    assert SOR = '1' report "Error in test case #493/2803" severity error;
    assert SOL = '0' report "Error in test case #493/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #494/2803" severity error;
    assert SOR = '1' report "Error in test case #494/2803" severity error;
    assert SOL = '0' report "Error in test case #494/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #495/2803" severity error;
    assert SOR = '1' report "Error in test case #495/2803" severity error;
    assert SOL = '0' report "Error in test case #495/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #496/2803" severity error;
    assert SOR = '1' report "Error in test case #496/2803" severity error;
    assert SOL = '0' report "Error in test case #496/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #497/2803" severity error;
    assert SOR = '1' report "Error in test case #497/2803" severity error;
    assert SOL = '0' report "Error in test case #497/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #498/2803" severity error;
    assert SOR = '1' report "Error in test case #498/2803" severity error;
    assert SOL = '0' report "Error in test case #498/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #499/2803" severity error;
    assert SOR = '1' report "Error in test case #499/2803" severity error;
    assert SOL = '0' report "Error in test case #499/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #500/2803" severity error;
    assert SOR = '1' report "Error in test case #500/2803" severity error;
    assert SOL = '0' report "Error in test case #500/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #501/2803" severity error;
    assert SOR = '1' report "Error in test case #501/2803" severity error;
    assert SOL = '0' report "Error in test case #501/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #502/2803" severity error;
    assert SOR = '1' report "Error in test case #502/2803" severity error;
    assert SOL = '0' report "Error in test case #502/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #503/2803" severity error;
    assert SOR = '1' report "Error in test case #503/2803" severity error;
    assert SOL = '0' report "Error in test case #503/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #504/2803" severity error;
    assert SOR = '1' report "Error in test case #504/2803" severity error;
    assert SOL = '0' report "Error in test case #504/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #505/2803" severity error;
    assert SOR = '1' report "Error in test case #505/2803" severity error;
    assert SOL = '0' report "Error in test case #505/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #506/2803" severity error;
    assert SOR = '1' report "Error in test case #506/2803" severity error;
    assert SOL = '0' report "Error in test case #506/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #507/2803" severity error;
    assert SOR = '1' report "Error in test case #507/2803" severity error;
    assert SOL = '0' report "Error in test case #507/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #508/2803" severity error;
    assert SOR = '1' report "Error in test case #508/2803" severity error;
    assert SOL = '0' report "Error in test case #508/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #509/2803" severity error;
    assert SOR = '1' report "Error in test case #509/2803" severity error;
    assert SOL = '0' report "Error in test case #509/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #510/2803" severity error;
    assert SOR = '1' report "Error in test case #510/2803" severity error;
    assert SOL = '0' report "Error in test case #510/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #511/2803" severity error;
    assert SOR = '1' report "Error in test case #511/2803" severity error;
    assert SOL = '0' report "Error in test case #511/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #512/2803" severity error;
    assert SOR = '1' report "Error in test case #512/2803" severity error;
    assert SOL = '0' report "Error in test case #512/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #513/2803" severity error;
    assert SOR = '1' report "Error in test case #513/2803" severity error;
    assert SOL = '0' report "Error in test case #513/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #514/2803" severity error;
    assert SOR = '1' report "Error in test case #514/2803" severity error;
    assert SOL = '0' report "Error in test case #514/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #515/2803" severity error;
    assert SOR = '1' report "Error in test case #515/2803" severity error;
    assert SOL = '0' report "Error in test case #515/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #516/2803" severity error;
    assert SOR = '1' report "Error in test case #516/2803" severity error;
    assert SOL = '0' report "Error in test case #516/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #517/2803" severity error;
    assert SOR = '1' report "Error in test case #517/2803" severity error;
    assert SOL = '0' report "Error in test case #517/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #518/2803" severity error;
    assert SOR = '1' report "Error in test case #518/2803" severity error;
    assert SOL = '0' report "Error in test case #518/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #519/2803" severity error;
    assert SOR = '1' report "Error in test case #519/2803" severity error;
    assert SOL = '0' report "Error in test case #519/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #520/2803" severity error;
    assert SOR = '1' report "Error in test case #520/2803" severity error;
    assert SOL = '0' report "Error in test case #520/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #521/2803" severity error;
    assert SOR = '1' report "Error in test case #521/2803" severity error;
    assert SOL = '0' report "Error in test case #521/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #522/2803" severity error;
    assert SOR = '1' report "Error in test case #522/2803" severity error;
    assert SOL = '0' report "Error in test case #522/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #523/2803" severity error;
    assert SOR = '1' report "Error in test case #523/2803" severity error;
    assert SOL = '0' report "Error in test case #523/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #524/2803" severity error;
    assert SOR = '1' report "Error in test case #524/2803" severity error;
    assert SOL = '0' report "Error in test case #524/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #525/2803" severity error;
    assert SOR = '1' report "Error in test case #525/2803" severity error;
    assert SOL = '0' report "Error in test case #525/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #526/2803" severity error;
    assert SOR = '1' report "Error in test case #526/2803" severity error;
    assert SOL = '1' report "Error in test case #526/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #527/2803" severity error;
    assert SOR = '1' report "Error in test case #527/2803" severity error;
    assert SOL = '1' report "Error in test case #527/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #528/2803" severity error;
    assert SOR = '1' report "Error in test case #528/2803" severity error;
    assert SOL = '1' report "Error in test case #528/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #529/2803" severity error;
    assert SOR = '1' report "Error in test case #529/2803" severity error;
    assert SOL = '1' report "Error in test case #529/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #530/2803" severity error;
    assert SOR = '1' report "Error in test case #530/2803" severity error;
    assert SOL = '1' report "Error in test case #530/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #531/2803" severity error;
    assert SOR = '1' report "Error in test case #531/2803" severity error;
    assert SOL = '1' report "Error in test case #531/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #532/2803" severity error;
    assert SOR = '1' report "Error in test case #532/2803" severity error;
    assert SOL = '1' report "Error in test case #532/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #533/2803" severity error;
    assert SOR = '1' report "Error in test case #533/2803" severity error;
    assert SOL = '1' report "Error in test case #533/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #534/2803" severity error;
    assert SOR = '1' report "Error in test case #534/2803" severity error;
    assert SOL = '1' report "Error in test case #534/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #535/2803" severity error;
    assert SOR = '1' report "Error in test case #535/2803" severity error;
    assert SOL = '1' report "Error in test case #535/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #536/2803" severity error;
    assert SOR = '1' report "Error in test case #536/2803" severity error;
    assert SOL = '0' report "Error in test case #536/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #537/2803" severity error;
    assert SOR = '1' report "Error in test case #537/2803" severity error;
    assert SOL = '0' report "Error in test case #537/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #538/2803" severity error;
    assert SOR = '1' report "Error in test case #538/2803" severity error;
    assert SOL = '0' report "Error in test case #538/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #539/2803" severity error;
    assert SOR = '1' report "Error in test case #539/2803" severity error;
    assert SOL = '0' report "Error in test case #539/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #540/2803" severity error;
    assert SOR = '1' report "Error in test case #540/2803" severity error;
    assert SOL = '0' report "Error in test case #540/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #541/2803" severity error;
    assert SOR = '1' report "Error in test case #541/2803" severity error;
    assert SOL = '0' report "Error in test case #541/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #542/2803" severity error;
    assert SOR = '1' report "Error in test case #542/2803" severity error;
    assert SOL = '0' report "Error in test case #542/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #543/2803" severity error;
    assert SOR = '1' report "Error in test case #543/2803" severity error;
    assert SOL = '0' report "Error in test case #543/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #544/2803" severity error;
    assert SOR = '1' report "Error in test case #544/2803" severity error;
    assert SOL = '1' report "Error in test case #544/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #545/2803" severity error;
    assert SOR = '1' report "Error in test case #545/2803" severity error;
    assert SOL = '1' report "Error in test case #545/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #546/2803" severity error;
    assert SOR = '1' report "Error in test case #546/2803" severity error;
    assert SOL = '1' report "Error in test case #546/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #547/2803" severity error;
    assert SOR = '1' report "Error in test case #547/2803" severity error;
    assert SOL = '1' report "Error in test case #547/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #548/2803" severity error;
    assert SOR = '1' report "Error in test case #548/2803" severity error;
    assert SOL = '1' report "Error in test case #548/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #549/2803" severity error;
    assert SOR = '1' report "Error in test case #549/2803" severity error;
    assert SOL = '1' report "Error in test case #549/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #550/2803" severity error;
    assert SOR = '1' report "Error in test case #550/2803" severity error;
    assert SOL = '1' report "Error in test case #550/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #551/2803" severity error;
    assert SOR = '1' report "Error in test case #551/2803" severity error;
    assert SOL = '1' report "Error in test case #551/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #552/2803" severity error;
    assert SOR = '1' report "Error in test case #552/2803" severity error;
    assert SOL = '1' report "Error in test case #552/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #553/2803" severity error;
    assert SOR = '1' report "Error in test case #553/2803" severity error;
    assert SOL = '1' report "Error in test case #553/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #554/2803" severity error;
    assert SOR = '1' report "Error in test case #554/2803" severity error;
    assert SOL = '1' report "Error in test case #554/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #555/2803" severity error;
    assert SOR = '1' report "Error in test case #555/2803" severity error;
    assert SOL = '1' report "Error in test case #555/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #556/2803" severity error;
    assert SOR = '1' report "Error in test case #556/2803" severity error;
    assert SOL = '1' report "Error in test case #556/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #557/2803" severity error;
    assert SOR = '1' report "Error in test case #557/2803" severity error;
    assert SOL = '1' report "Error in test case #557/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #558/2803" severity error;
    assert SOR = '1' report "Error in test case #558/2803" severity error;
    assert SOL = '1' report "Error in test case #558/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #559/2803" severity error;
    assert SOR = '1' report "Error in test case #559/2803" severity error;
    assert SOL = '1' report "Error in test case #559/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #560/2803" severity error;
    assert SOR = '1' report "Error in test case #560/2803" severity error;
    assert SOL = '1' report "Error in test case #560/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #561/2803" severity error;
    assert SOR = '1' report "Error in test case #561/2803" severity error;
    assert SOL = '1' report "Error in test case #561/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #562/2803" severity error;
    assert SOR = '1' report "Error in test case #562/2803" severity error;
    assert SOL = '1' report "Error in test case #562/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #563/2803" severity error;
    assert SOR = '1' report "Error in test case #563/2803" severity error;
    assert SOL = '1' report "Error in test case #563/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #564/2803" severity error;
    assert SOR = '1' report "Error in test case #564/2803" severity error;
    assert SOL = '1' report "Error in test case #564/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #565/2803" severity error;
    assert SOR = '1' report "Error in test case #565/2803" severity error;
    assert SOL = '1' report "Error in test case #565/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #566/2803" severity error;
    assert SOR = '1' report "Error in test case #566/2803" severity error;
    assert SOL = '1' report "Error in test case #566/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #567/2803" severity error;
    assert SOR = '1' report "Error in test case #567/2803" severity error;
    assert SOL = '1' report "Error in test case #567/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #568/2803" severity error;
    assert SOR = '1' report "Error in test case #568/2803" severity error;
    assert SOL = '1' report "Error in test case #568/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #569/2803" severity error;
    assert SOR = '1' report "Error in test case #569/2803" severity error;
    assert SOL = '1' report "Error in test case #569/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #570/2803" severity error;
    assert SOR = '1' report "Error in test case #570/2803" severity error;
    assert SOL = '1' report "Error in test case #570/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #571/2803" severity error;
    assert SOR = '1' report "Error in test case #571/2803" severity error;
    assert SOL = '1' report "Error in test case #571/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #572/2803" severity error;
    assert SOR = '1' report "Error in test case #572/2803" severity error;
    assert SOL = '1' report "Error in test case #572/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #573/2803" severity error;
    assert SOR = '1' report "Error in test case #573/2803" severity error;
    assert SOL = '1' report "Error in test case #573/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #574/2803" severity error;
    assert SOR = '1' report "Error in test case #574/2803" severity error;
    assert SOL = '1' report "Error in test case #574/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #575/2803" severity error;
    assert SOR = '1' report "Error in test case #575/2803" severity error;
    assert SOL = '1' report "Error in test case #575/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #576/2803" severity error;
    assert SOR = '1' report "Error in test case #576/2803" severity error;
    assert SOL = '0' report "Error in test case #576/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #577/2803" severity error;
    assert SOR = '1' report "Error in test case #577/2803" severity error;
    assert SOL = '0' report "Error in test case #577/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #578/2803" severity error;
    assert SOR = '1' report "Error in test case #578/2803" severity error;
    assert SOL = '0' report "Error in test case #578/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #579/2803" severity error;
    assert SOR = '1' report "Error in test case #579/2803" severity error;
    assert SOL = '0' report "Error in test case #579/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #580/2803" severity error;
    assert SOR = '1' report "Error in test case #580/2803" severity error;
    assert SOL = '0' report "Error in test case #580/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #581/2803" severity error;
    assert SOR = '1' report "Error in test case #581/2803" severity error;
    assert SOL = '0' report "Error in test case #581/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #582/2803" severity error;
    assert SOR = '1' report "Error in test case #582/2803" severity error;
    assert SOL = '0' report "Error in test case #582/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #583/2803" severity error;
    assert SOR = '1' report "Error in test case #583/2803" severity error;
    assert SOL = '0' report "Error in test case #583/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #584/2803" severity error;
    assert SOR = '1' report "Error in test case #584/2803" severity error;
    assert SOL = '0' report "Error in test case #584/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #585/2803" severity error;
    assert SOR = '1' report "Error in test case #585/2803" severity error;
    assert SOL = '0' report "Error in test case #585/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #586/2803" severity error;
    assert SOR = '1' report "Error in test case #586/2803" severity error;
    assert SOL = '0' report "Error in test case #586/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #587/2803" severity error;
    assert SOR = '1' report "Error in test case #587/2803" severity error;
    assert SOL = '0' report "Error in test case #587/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #588/2803" severity error;
    assert SOR = '1' report "Error in test case #588/2803" severity error;
    assert SOL = '0' report "Error in test case #588/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #589/2803" severity error;
    assert SOR = '1' report "Error in test case #589/2803" severity error;
    assert SOL = '0' report "Error in test case #589/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #590/2803" severity error;
    assert SOR = '1' report "Error in test case #590/2803" severity error;
    assert SOL = '0' report "Error in test case #590/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #591/2803" severity error;
    assert SOR = '1' report "Error in test case #591/2803" severity error;
    assert SOL = '0' report "Error in test case #591/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #592/2803" severity error;
    assert SOR = '1' report "Error in test case #592/2803" severity error;
    assert SOL = '0' report "Error in test case #592/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #593/2803" severity error;
    assert SOR = '1' report "Error in test case #593/2803" severity error;
    assert SOL = '0' report "Error in test case #593/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #594/2803" severity error;
    assert SOR = '1' report "Error in test case #594/2803" severity error;
    assert SOL = '0' report "Error in test case #594/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #595/2803" severity error;
    assert SOR = '1' report "Error in test case #595/2803" severity error;
    assert SOL = '0' report "Error in test case #595/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #596/2803" severity error;
    assert SOR = '1' report "Error in test case #596/2803" severity error;
    assert SOL = '0' report "Error in test case #596/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #597/2803" severity error;
    assert SOR = '1' report "Error in test case #597/2803" severity error;
    assert SOL = '0' report "Error in test case #597/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #598/2803" severity error;
    assert SOR = '1' report "Error in test case #598/2803" severity error;
    assert SOL = '0' report "Error in test case #598/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #599/2803" severity error;
    assert SOR = '1' report "Error in test case #599/2803" severity error;
    assert SOL = '0' report "Error in test case #599/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #600/2803" severity error;
    assert SOR = '1' report "Error in test case #600/2803" severity error;
    assert SOL = '0' report "Error in test case #600/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #601/2803" severity error;
    assert SOR = '1' report "Error in test case #601/2803" severity error;
    assert SOL = '0' report "Error in test case #601/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #602/2803" severity error;
    assert SOR = '1' report "Error in test case #602/2803" severity error;
    assert SOL = '0' report "Error in test case #602/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #603/2803" severity error;
    assert SOR = '0' report "Error in test case #603/2803" severity error;
    assert SOL = '0' report "Error in test case #603/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #604/2803" severity error;
    assert SOR = '0' report "Error in test case #604/2803" severity error;
    assert SOL = '0' report "Error in test case #604/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #605/2803" severity error;
    assert SOR = '0' report "Error in test case #605/2803" severity error;
    assert SOL = '0' report "Error in test case #605/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #606/2803" severity error;
    assert SOR = '0' report "Error in test case #606/2803" severity error;
    assert SOL = '0' report "Error in test case #606/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #607/2803" severity error;
    assert SOR = '0' report "Error in test case #607/2803" severity error;
    assert SOL = '0' report "Error in test case #607/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #608/2803" severity error;
    assert SOR = '0' report "Error in test case #608/2803" severity error;
    assert SOL = '0' report "Error in test case #608/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #609/2803" severity error;
    assert SOR = '0' report "Error in test case #609/2803" severity error;
    assert SOL = '0' report "Error in test case #609/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #610/2803" severity error;
    assert SOR = '0' report "Error in test case #610/2803" severity error;
    assert SOL = '0' report "Error in test case #610/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #611/2803" severity error;
    assert SOR = '0' report "Error in test case #611/2803" severity error;
    assert SOL = '0' report "Error in test case #611/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #612/2803" severity error;
    assert SOR = '0' report "Error in test case #612/2803" severity error;
    assert SOL = '0' report "Error in test case #612/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #613/2803" severity error;
    assert SOR = '0' report "Error in test case #613/2803" severity error;
    assert SOL = '0' report "Error in test case #613/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #614/2803" severity error;
    assert SOR = '0' report "Error in test case #614/2803" severity error;
    assert SOL = '0' report "Error in test case #614/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #615/2803" severity error;
    assert SOR = '0' report "Error in test case #615/2803" severity error;
    assert SOL = '0' report "Error in test case #615/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #616/2803" severity error;
    assert SOR = '0' report "Error in test case #616/2803" severity error;
    assert SOL = '0' report "Error in test case #616/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #617/2803" severity error;
    assert SOR = '0' report "Error in test case #617/2803" severity error;
    assert SOL = '0' report "Error in test case #617/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #618/2803" severity error;
    assert SOR = '0' report "Error in test case #618/2803" severity error;
    assert SOL = '0' report "Error in test case #618/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #619/2803" severity error;
    assert SOR = '0' report "Error in test case #619/2803" severity error;
    assert SOL = '0' report "Error in test case #619/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #620/2803" severity error;
    assert SOR = '0' report "Error in test case #620/2803" severity error;
    assert SOL = '0' report "Error in test case #620/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #621/2803" severity error;
    assert SOR = '0' report "Error in test case #621/2803" severity error;
    assert SOL = '0' report "Error in test case #621/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #622/2803" severity error;
    assert SOR = '0' report "Error in test case #622/2803" severity error;
    assert SOL = '0' report "Error in test case #622/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #623/2803" severity error;
    assert SOR = '0' report "Error in test case #623/2803" severity error;
    assert SOL = '0' report "Error in test case #623/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #624/2803" severity error;
    assert SOR = '0' report "Error in test case #624/2803" severity error;
    assert SOL = '1' report "Error in test case #624/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #625/2803" severity error;
    assert SOR = '0' report "Error in test case #625/2803" severity error;
    assert SOL = '1' report "Error in test case #625/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #626/2803" severity error;
    assert SOR = '0' report "Error in test case #626/2803" severity error;
    assert SOL = '1' report "Error in test case #626/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #627/2803" severity error;
    assert SOR = '0' report "Error in test case #627/2803" severity error;
    assert SOL = '1' report "Error in test case #627/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #628/2803" severity error;
    assert SOR = '0' report "Error in test case #628/2803" severity error;
    assert SOL = '1' report "Error in test case #628/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #629/2803" severity error;
    assert SOR = '1' report "Error in test case #629/2803" severity error;
    assert SOL = '1' report "Error in test case #629/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #630/2803" severity error;
    assert SOR = '1' report "Error in test case #630/2803" severity error;
    assert SOL = '1' report "Error in test case #630/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #631/2803" severity error;
    assert SOR = '1' report "Error in test case #631/2803" severity error;
    assert SOL = '1' report "Error in test case #631/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #632/2803" severity error;
    assert SOR = '1' report "Error in test case #632/2803" severity error;
    assert SOL = '0' report "Error in test case #632/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #633/2803" severity error;
    assert SOR = '1' report "Error in test case #633/2803" severity error;
    assert SOL = '0' report "Error in test case #633/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #634/2803" severity error;
    assert SOR = '1' report "Error in test case #634/2803" severity error;
    assert SOL = '0' report "Error in test case #634/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #635/2803" severity error;
    assert SOR = '1' report "Error in test case #635/2803" severity error;
    assert SOL = '0' report "Error in test case #635/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #636/2803" severity error;
    assert SOR = '1' report "Error in test case #636/2803" severity error;
    assert SOL = '0' report "Error in test case #636/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #637/2803" severity error;
    assert SOR = '1' report "Error in test case #637/2803" severity error;
    assert SOL = '0' report "Error in test case #637/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #638/2803" severity error;
    assert SOR = '1' report "Error in test case #638/2803" severity error;
    assert SOL = '0' report "Error in test case #638/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #639/2803" severity error;
    assert SOR = '1' report "Error in test case #639/2803" severity error;
    assert SOL = '0' report "Error in test case #639/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #640/2803" severity error;
    assert SOR = '1' report "Error in test case #640/2803" severity error;
    assert SOL = '0' report "Error in test case #640/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #641/2803" severity error;
    assert SOR = '1' report "Error in test case #641/2803" severity error;
    assert SOL = '0' report "Error in test case #641/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #642/2803" severity error;
    assert SOR = '1' report "Error in test case #642/2803" severity error;
    assert SOL = '0' report "Error in test case #642/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #643/2803" severity error;
    assert SOR = '1' report "Error in test case #643/2803" severity error;
    assert SOL = '0' report "Error in test case #643/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #644/2803" severity error;
    assert SOR = '1' report "Error in test case #644/2803" severity error;
    assert SOL = '0' report "Error in test case #644/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #645/2803" severity error;
    assert SOR = '1' report "Error in test case #645/2803" severity error;
    assert SOL = '0' report "Error in test case #645/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #646/2803" severity error;
    assert SOR = '1' report "Error in test case #646/2803" severity error;
    assert SOL = '0' report "Error in test case #646/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #647/2803" severity error;
    assert SOR = '1' report "Error in test case #647/2803" severity error;
    assert SOL = '0' report "Error in test case #647/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10011111" report "Error in test case #648/2803" severity error;
    assert SOR = '1' report "Error in test case #648/2803" severity error;
    assert SOL = '1' report "Error in test case #648/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10011111" report "Error in test case #649/2803" severity error;
    assert SOR = '1' report "Error in test case #649/2803" severity error;
    assert SOL = '1' report "Error in test case #649/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #650/2803" severity error;
    assert SOR = '0' report "Error in test case #650/2803" severity error;
    assert SOL = '0' report "Error in test case #650/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #651/2803" severity error;
    assert SOR = '0' report "Error in test case #651/2803" severity error;
    assert SOL = '0' report "Error in test case #651/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #652/2803" severity error;
    assert SOR = '0' report "Error in test case #652/2803" severity error;
    assert SOL = '0' report "Error in test case #652/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #653/2803" severity error;
    assert SOR = '0' report "Error in test case #653/2803" severity error;
    assert SOL = '0' report "Error in test case #653/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #654/2803" severity error;
    assert SOR = '0' report "Error in test case #654/2803" severity error;
    assert SOL = '0' report "Error in test case #654/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #655/2803" severity error;
    assert SOR = '0' report "Error in test case #655/2803" severity error;
    assert SOL = '0' report "Error in test case #655/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #656/2803" severity error;
    assert SOR = '0' report "Error in test case #656/2803" severity error;
    assert SOL = '0' report "Error in test case #656/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #657/2803" severity error;
    assert SOR = '0' report "Error in test case #657/2803" severity error;
    assert SOL = '0' report "Error in test case #657/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #658/2803" severity error;
    assert SOR = '0' report "Error in test case #658/2803" severity error;
    assert SOL = '0' report "Error in test case #658/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #659/2803" severity error;
    assert SOR = '0' report "Error in test case #659/2803" severity error;
    assert SOL = '0' report "Error in test case #659/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #660/2803" severity error;
    assert SOR = '0' report "Error in test case #660/2803" severity error;
    assert SOL = '0' report "Error in test case #660/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #661/2803" severity error;
    assert SOR = '0' report "Error in test case #661/2803" severity error;
    assert SOL = '0' report "Error in test case #661/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #662/2803" severity error;
    assert SOR = '0' report "Error in test case #662/2803" severity error;
    assert SOL = '0' report "Error in test case #662/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #663/2803" severity error;
    assert SOR = '0' report "Error in test case #663/2803" severity error;
    assert SOL = '0' report "Error in test case #663/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #664/2803" severity error;
    assert SOR = '0' report "Error in test case #664/2803" severity error;
    assert SOL = '1' report "Error in test case #664/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #665/2803" severity error;
    assert SOR = '0' report "Error in test case #665/2803" severity error;
    assert SOL = '1' report "Error in test case #665/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #666/2803" severity error;
    assert SOR = '0' report "Error in test case #666/2803" severity error;
    assert SOL = '1' report "Error in test case #666/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #667/2803" severity error;
    assert SOR = '0' report "Error in test case #667/2803" severity error;
    assert SOL = '1' report "Error in test case #667/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #668/2803" severity error;
    assert SOR = '0' report "Error in test case #668/2803" severity error;
    assert SOL = '1' report "Error in test case #668/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #669/2803" severity error;
    assert SOR = '0' report "Error in test case #669/2803" severity error;
    assert SOL = '1' report "Error in test case #669/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #670/2803" severity error;
    assert SOR = '0' report "Error in test case #670/2803" severity error;
    assert SOL = '1' report "Error in test case #670/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10000000" report "Error in test case #671/2803" severity error;
    assert SOR = '0' report "Error in test case #671/2803" severity error;
    assert SOL = '1' report "Error in test case #671/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11000000" report "Error in test case #672/2803" severity error;
    assert SOR = '0' report "Error in test case #672/2803" severity error;
    assert SOL = '1' report "Error in test case #672/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11000000" report "Error in test case #673/2803" severity error;
    assert SOR = '0' report "Error in test case #673/2803" severity error;
    assert SOL = '1' report "Error in test case #673/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11000000" report "Error in test case #674/2803" severity error;
    assert SOR = '0' report "Error in test case #674/2803" severity error;
    assert SOL = '1' report "Error in test case #674/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11000000" report "Error in test case #675/2803" severity error;
    assert SOR = '0' report "Error in test case #675/2803" severity error;
    assert SOL = '1' report "Error in test case #675/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11000000" report "Error in test case #676/2803" severity error;
    assert SOR = '0' report "Error in test case #676/2803" severity error;
    assert SOL = '1' report "Error in test case #676/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11000000" report "Error in test case #677/2803" severity error;
    assert SOR = '0' report "Error in test case #677/2803" severity error;
    assert SOL = '1' report "Error in test case #677/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11000000" report "Error in test case #678/2803" severity error;
    assert SOR = '0' report "Error in test case #678/2803" severity error;
    assert SOL = '1' report "Error in test case #678/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11000000" report "Error in test case #679/2803" severity error;
    assert SOR = '0' report "Error in test case #679/2803" severity error;
    assert SOL = '1' report "Error in test case #679/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01100000" report "Error in test case #680/2803" severity error;
    assert SOR = '0' report "Error in test case #680/2803" severity error;
    assert SOL = '0' report "Error in test case #680/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01100000" report "Error in test case #681/2803" severity error;
    assert SOR = '0' report "Error in test case #681/2803" severity error;
    assert SOL = '0' report "Error in test case #681/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01100000" report "Error in test case #682/2803" severity error;
    assert SOR = '0' report "Error in test case #682/2803" severity error;
    assert SOL = '0' report "Error in test case #682/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01100000" report "Error in test case #683/2803" severity error;
    assert SOR = '0' report "Error in test case #683/2803" severity error;
    assert SOL = '0' report "Error in test case #683/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01100000" report "Error in test case #684/2803" severity error;
    assert SOR = '0' report "Error in test case #684/2803" severity error;
    assert SOL = '0' report "Error in test case #684/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01100000" report "Error in test case #685/2803" severity error;
    assert SOR = '0' report "Error in test case #685/2803" severity error;
    assert SOL = '0' report "Error in test case #685/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01100000" report "Error in test case #686/2803" severity error;
    assert SOR = '0' report "Error in test case #686/2803" severity error;
    assert SOL = '0' report "Error in test case #686/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01100000" report "Error in test case #687/2803" severity error;
    assert SOR = '0' report "Error in test case #687/2803" severity error;
    assert SOL = '0' report "Error in test case #687/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10110000" report "Error in test case #688/2803" severity error;
    assert SOR = '0' report "Error in test case #688/2803" severity error;
    assert SOL = '1' report "Error in test case #688/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10110000" report "Error in test case #689/2803" severity error;
    assert SOR = '0' report "Error in test case #689/2803" severity error;
    assert SOL = '1' report "Error in test case #689/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10110000" report "Error in test case #690/2803" severity error;
    assert SOR = '0' report "Error in test case #690/2803" severity error;
    assert SOL = '1' report "Error in test case #690/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10110000" report "Error in test case #691/2803" severity error;
    assert SOR = '0' report "Error in test case #691/2803" severity error;
    assert SOL = '1' report "Error in test case #691/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10110000" report "Error in test case #692/2803" severity error;
    assert SOR = '0' report "Error in test case #692/2803" severity error;
    assert SOL = '1' report "Error in test case #692/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10110000" report "Error in test case #693/2803" severity error;
    assert SOR = '0' report "Error in test case #693/2803" severity error;
    assert SOL = '1' report "Error in test case #693/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10110000" report "Error in test case #694/2803" severity error;
    assert SOR = '0' report "Error in test case #694/2803" severity error;
    assert SOL = '1' report "Error in test case #694/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10110000" report "Error in test case #695/2803" severity error;
    assert SOR = '0' report "Error in test case #695/2803" severity error;
    assert SOL = '1' report "Error in test case #695/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01011000" report "Error in test case #696/2803" severity error;
    assert SOR = '0' report "Error in test case #696/2803" severity error;
    assert SOL = '0' report "Error in test case #696/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01011000" report "Error in test case #697/2803" severity error;
    assert SOR = '0' report "Error in test case #697/2803" severity error;
    assert SOL = '0' report "Error in test case #697/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01011000" report "Error in test case #698/2803" severity error;
    assert SOR = '0' report "Error in test case #698/2803" severity error;
    assert SOL = '0' report "Error in test case #698/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01011000" report "Error in test case #699/2803" severity error;
    assert SOR = '0' report "Error in test case #699/2803" severity error;
    assert SOL = '0' report "Error in test case #699/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01011000" report "Error in test case #700/2803" severity error;
    assert SOR = '0' report "Error in test case #700/2803" severity error;
    assert SOL = '0' report "Error in test case #700/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01011000" report "Error in test case #701/2803" severity error;
    assert SOR = '0' report "Error in test case #701/2803" severity error;
    assert SOL = '0' report "Error in test case #701/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01011000" report "Error in test case #702/2803" severity error;
    assert SOR = '0' report "Error in test case #702/2803" severity error;
    assert SOL = '0' report "Error in test case #702/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01011000" report "Error in test case #703/2803" severity error;
    assert SOR = '0' report "Error in test case #703/2803" severity error;
    assert SOL = '0' report "Error in test case #703/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10101100" report "Error in test case #704/2803" severity error;
    assert SOR = '0' report "Error in test case #704/2803" severity error;
    assert SOL = '1' report "Error in test case #704/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10101100" report "Error in test case #705/2803" severity error;
    assert SOR = '0' report "Error in test case #705/2803" severity error;
    assert SOL = '1' report "Error in test case #705/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10101100" report "Error in test case #706/2803" severity error;
    assert SOR = '0' report "Error in test case #706/2803" severity error;
    assert SOL = '1' report "Error in test case #706/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10101100" report "Error in test case #707/2803" severity error;
    assert SOR = '0' report "Error in test case #707/2803" severity error;
    assert SOL = '1' report "Error in test case #707/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10101100" report "Error in test case #708/2803" severity error;
    assert SOR = '0' report "Error in test case #708/2803" severity error;
    assert SOL = '1' report "Error in test case #708/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10101100" report "Error in test case #709/2803" severity error;
    assert SOR = '0' report "Error in test case #709/2803" severity error;
    assert SOL = '1' report "Error in test case #709/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10101100" report "Error in test case #710/2803" severity error;
    assert SOR = '0' report "Error in test case #710/2803" severity error;
    assert SOL = '1' report "Error in test case #710/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10101100" report "Error in test case #711/2803" severity error;
    assert SOR = '0' report "Error in test case #711/2803" severity error;
    assert SOL = '1' report "Error in test case #711/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01010110" report "Error in test case #712/2803" severity error;
    assert SOR = '0' report "Error in test case #712/2803" severity error;
    assert SOL = '0' report "Error in test case #712/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01010110" report "Error in test case #713/2803" severity error;
    assert SOR = '0' report "Error in test case #713/2803" severity error;
    assert SOL = '0' report "Error in test case #713/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01010110" report "Error in test case #714/2803" severity error;
    assert SOR = '0' report "Error in test case #714/2803" severity error;
    assert SOL = '0' report "Error in test case #714/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01010110" report "Error in test case #715/2803" severity error;
    assert SOR = '0' report "Error in test case #715/2803" severity error;
    assert SOL = '0' report "Error in test case #715/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01010110" report "Error in test case #716/2803" severity error;
    assert SOR = '0' report "Error in test case #716/2803" severity error;
    assert SOL = '0' report "Error in test case #716/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01010110" report "Error in test case #717/2803" severity error;
    assert SOR = '0' report "Error in test case #717/2803" severity error;
    assert SOL = '0' report "Error in test case #717/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01010110" report "Error in test case #718/2803" severity error;
    assert SOR = '0' report "Error in test case #718/2803" severity error;
    assert SOL = '0' report "Error in test case #718/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01010110" report "Error in test case #719/2803" severity error;
    assert SOR = '0' report "Error in test case #719/2803" severity error;
    assert SOL = '0' report "Error in test case #719/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #720/2803" severity error;
    assert SOR = '1' report "Error in test case #720/2803" severity error;
    assert SOL = '1' report "Error in test case #720/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #721/2803" severity error;
    assert SOR = '1' report "Error in test case #721/2803" severity error;
    assert SOL = '1' report "Error in test case #721/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #722/2803" severity error;
    assert SOR = '1' report "Error in test case #722/2803" severity error;
    assert SOL = '1' report "Error in test case #722/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #723/2803" severity error;
    assert SOR = '1' report "Error in test case #723/2803" severity error;
    assert SOL = '1' report "Error in test case #723/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #724/2803" severity error;
    assert SOR = '1' report "Error in test case #724/2803" severity error;
    assert SOL = '1' report "Error in test case #724/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #725/2803" severity error;
    assert SOR = '1' report "Error in test case #725/2803" severity error;
    assert SOL = '1' report "Error in test case #725/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #726/2803" severity error;
    assert SOR = '1' report "Error in test case #726/2803" severity error;
    assert SOL = '1' report "Error in test case #726/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #727/2803" severity error;
    assert SOR = '1' report "Error in test case #727/2803" severity error;
    assert SOL = '1' report "Error in test case #727/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #728/2803" severity error;
    assert SOR = '1' report "Error in test case #728/2803" severity error;
    assert SOL = '1' report "Error in test case #728/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #729/2803" severity error;
    assert SOR = '1' report "Error in test case #729/2803" severity error;
    assert SOL = '1' report "Error in test case #729/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #730/2803" severity error;
    assert SOR = '1' report "Error in test case #730/2803" severity error;
    assert SOL = '1' report "Error in test case #730/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #731/2803" severity error;
    assert SOR = '1' report "Error in test case #731/2803" severity error;
    assert SOL = '1' report "Error in test case #731/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #732/2803" severity error;
    assert SOR = '1' report "Error in test case #732/2803" severity error;
    assert SOL = '1' report "Error in test case #732/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #733/2803" severity error;
    assert SOR = '1' report "Error in test case #733/2803" severity error;
    assert SOL = '1' report "Error in test case #733/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #734/2803" severity error;
    assert SOR = '1' report "Error in test case #734/2803" severity error;
    assert SOL = '1' report "Error in test case #734/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #735/2803" severity error;
    assert SOR = '1' report "Error in test case #735/2803" severity error;
    assert SOL = '1' report "Error in test case #735/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #736/2803" severity error;
    assert SOR = '1' report "Error in test case #736/2803" severity error;
    assert SOL = '0' report "Error in test case #736/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #737/2803" severity error;
    assert SOR = '1' report "Error in test case #737/2803" severity error;
    assert SOL = '0' report "Error in test case #737/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #738/2803" severity error;
    assert SOR = '1' report "Error in test case #738/2803" severity error;
    assert SOL = '0' report "Error in test case #738/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #739/2803" severity error;
    assert SOR = '1' report "Error in test case #739/2803" severity error;
    assert SOL = '0' report "Error in test case #739/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #740/2803" severity error;
    assert SOR = '1' report "Error in test case #740/2803" severity error;
    assert SOL = '0' report "Error in test case #740/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #741/2803" severity error;
    assert SOR = '1' report "Error in test case #741/2803" severity error;
    assert SOL = '0' report "Error in test case #741/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #742/2803" severity error;
    assert SOR = '1' report "Error in test case #742/2803" severity error;
    assert SOL = '0' report "Error in test case #742/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #743/2803" severity error;
    assert SOR = '1' report "Error in test case #743/2803" severity error;
    assert SOL = '0' report "Error in test case #743/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #744/2803" severity error;
    assert SOR = '1' report "Error in test case #744/2803" severity error;
    assert SOL = '1' report "Error in test case #744/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #745/2803" severity error;
    assert SOR = '1' report "Error in test case #745/2803" severity error;
    assert SOL = '1' report "Error in test case #745/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #746/2803" severity error;
    assert SOR = '1' report "Error in test case #746/2803" severity error;
    assert SOL = '1' report "Error in test case #746/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #747/2803" severity error;
    assert SOR = '1' report "Error in test case #747/2803" severity error;
    assert SOL = '1' report "Error in test case #747/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #748/2803" severity error;
    assert SOR = '1' report "Error in test case #748/2803" severity error;
    assert SOL = '1' report "Error in test case #748/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #749/2803" severity error;
    assert SOR = '1' report "Error in test case #749/2803" severity error;
    assert SOL = '1' report "Error in test case #749/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #750/2803" severity error;
    assert SOR = '1' report "Error in test case #750/2803" severity error;
    assert SOL = '1' report "Error in test case #750/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10111111" report "Error in test case #751/2803" severity error;
    assert SOR = '1' report "Error in test case #751/2803" severity error;
    assert SOL = '1' report "Error in test case #751/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01011111" report "Error in test case #752/2803" severity error;
    assert SOR = '1' report "Error in test case #752/2803" severity error;
    assert SOL = '0' report "Error in test case #752/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01011111" report "Error in test case #753/2803" severity error;
    assert SOR = '1' report "Error in test case #753/2803" severity error;
    assert SOL = '0' report "Error in test case #753/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01011111" report "Error in test case #754/2803" severity error;
    assert SOR = '1' report "Error in test case #754/2803" severity error;
    assert SOL = '0' report "Error in test case #754/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01011111" report "Error in test case #755/2803" severity error;
    assert SOR = '1' report "Error in test case #755/2803" severity error;
    assert SOL = '0' report "Error in test case #755/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01011111" report "Error in test case #756/2803" severity error;
    assert SOR = '1' report "Error in test case #756/2803" severity error;
    assert SOL = '0' report "Error in test case #756/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01011111" report "Error in test case #757/2803" severity error;
    assert SOR = '1' report "Error in test case #757/2803" severity error;
    assert SOL = '0' report "Error in test case #757/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01011111" report "Error in test case #758/2803" severity error;
    assert SOR = '1' report "Error in test case #758/2803" severity error;
    assert SOL = '0' report "Error in test case #758/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01011111" report "Error in test case #759/2803" severity error;
    assert SOR = '1' report "Error in test case #759/2803" severity error;
    assert SOL = '0' report "Error in test case #759/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00101111" report "Error in test case #760/2803" severity error;
    assert SOR = '1' report "Error in test case #760/2803" severity error;
    assert SOL = '0' report "Error in test case #760/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00101111" report "Error in test case #761/2803" severity error;
    assert SOR = '1' report "Error in test case #761/2803" severity error;
    assert SOL = '0' report "Error in test case #761/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00101111" report "Error in test case #762/2803" severity error;
    assert SOR = '1' report "Error in test case #762/2803" severity error;
    assert SOL = '0' report "Error in test case #762/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00101111" report "Error in test case #763/2803" severity error;
    assert SOR = '1' report "Error in test case #763/2803" severity error;
    assert SOL = '0' report "Error in test case #763/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00101111" report "Error in test case #764/2803" severity error;
    assert SOR = '1' report "Error in test case #764/2803" severity error;
    assert SOL = '0' report "Error in test case #764/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00101111" report "Error in test case #765/2803" severity error;
    assert SOR = '1' report "Error in test case #765/2803" severity error;
    assert SOL = '0' report "Error in test case #765/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00101111" report "Error in test case #766/2803" severity error;
    assert SOR = '1' report "Error in test case #766/2803" severity error;
    assert SOL = '0' report "Error in test case #766/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00101111" report "Error in test case #767/2803" severity error;
    assert SOR = '1' report "Error in test case #767/2803" severity error;
    assert SOL = '0' report "Error in test case #767/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010111" report "Error in test case #768/2803" severity error;
    assert SOR = '1' report "Error in test case #768/2803" severity error;
    assert SOL = '1' report "Error in test case #768/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "10010111" report "Error in test case #769/2803" severity error;
    assert SOR = '1' report "Error in test case #769/2803" severity error;
    assert SOL = '1' report "Error in test case #769/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10010111" report "Error in test case #770/2803" severity error;
    assert SOR = '1' report "Error in test case #770/2803" severity error;
    assert SOL = '1' report "Error in test case #770/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10010111" report "Error in test case #771/2803" severity error;
    assert SOR = '1' report "Error in test case #771/2803" severity error;
    assert SOL = '1' report "Error in test case #771/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10010111" report "Error in test case #772/2803" severity error;
    assert SOR = '1' report "Error in test case #772/2803" severity error;
    assert SOL = '1' report "Error in test case #772/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10010111" report "Error in test case #773/2803" severity error;
    assert SOR = '1' report "Error in test case #773/2803" severity error;
    assert SOL = '1' report "Error in test case #773/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10010111" report "Error in test case #774/2803" severity error;
    assert SOR = '1' report "Error in test case #774/2803" severity error;
    assert SOL = '1' report "Error in test case #774/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "10010111" report "Error in test case #775/2803" severity error;
    assert SOR = '1' report "Error in test case #775/2803" severity error;
    assert SOL = '1' report "Error in test case #775/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01001011" report "Error in test case #776/2803" severity error;
    assert SOR = '1' report "Error in test case #776/2803" severity error;
    assert SOL = '0' report "Error in test case #776/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01001011" report "Error in test case #777/2803" severity error;
    assert SOR = '1' report "Error in test case #777/2803" severity error;
    assert SOL = '0' report "Error in test case #777/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #778/2803" severity error;
    assert SOR = '1' report "Error in test case #778/2803" severity error;
    assert SOL = '1' report "Error in test case #778/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #779/2803" severity error;
    assert SOR = '1' report "Error in test case #779/2803" severity error;
    assert SOL = '1' report "Error in test case #779/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #780/2803" severity error;
    assert SOR = '1' report "Error in test case #780/2803" severity error;
    assert SOL = '1' report "Error in test case #780/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #781/2803" severity error;
    assert SOR = '1' report "Error in test case #781/2803" severity error;
    assert SOL = '1' report "Error in test case #781/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #782/2803" severity error;
    assert SOR = '1' report "Error in test case #782/2803" severity error;
    assert SOL = '1' report "Error in test case #782/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #783/2803" severity error;
    assert SOR = '1' report "Error in test case #783/2803" severity error;
    assert SOL = '1' report "Error in test case #783/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #784/2803" severity error;
    assert SOR = '1' report "Error in test case #784/2803" severity error;
    assert SOL = '1' report "Error in test case #784/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #785/2803" severity error;
    assert SOR = '1' report "Error in test case #785/2803" severity error;
    assert SOL = '1' report "Error in test case #785/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #786/2803" severity error;
    assert SOR = '1' report "Error in test case #786/2803" severity error;
    assert SOL = '1' report "Error in test case #786/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #787/2803" severity error;
    assert SOR = '1' report "Error in test case #787/2803" severity error;
    assert SOL = '1' report "Error in test case #787/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #788/2803" severity error;
    assert SOR = '1' report "Error in test case #788/2803" severity error;
    assert SOL = '1' report "Error in test case #788/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #789/2803" severity error;
    assert SOR = '1' report "Error in test case #789/2803" severity error;
    assert SOL = '1' report "Error in test case #789/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #790/2803" severity error;
    assert SOR = '1' report "Error in test case #790/2803" severity error;
    assert SOL = '1' report "Error in test case #790/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #791/2803" severity error;
    assert SOR = '1' report "Error in test case #791/2803" severity error;
    assert SOL = '1' report "Error in test case #791/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #792/2803" severity error;
    assert SOR = '1' report "Error in test case #792/2803" severity error;
    assert SOL = '0' report "Error in test case #792/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #793/2803" severity error;
    assert SOR = '1' report "Error in test case #793/2803" severity error;
    assert SOL = '0' report "Error in test case #793/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #794/2803" severity error;
    assert SOR = '1' report "Error in test case #794/2803" severity error;
    assert SOL = '0' report "Error in test case #794/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #795/2803" severity error;
    assert SOR = '1' report "Error in test case #795/2803" severity error;
    assert SOL = '0' report "Error in test case #795/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #796/2803" severity error;
    assert SOR = '1' report "Error in test case #796/2803" severity error;
    assert SOL = '1' report "Error in test case #796/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #797/2803" severity error;
    assert SOR = '1' report "Error in test case #797/2803" severity error;
    assert SOL = '1' report "Error in test case #797/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #798/2803" severity error;
    assert SOR = '1' report "Error in test case #798/2803" severity error;
    assert SOL = '1' report "Error in test case #798/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #799/2803" severity error;
    assert SOR = '1' report "Error in test case #799/2803" severity error;
    assert SOL = '1' report "Error in test case #799/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #800/2803" severity error;
    assert SOR = '1' report "Error in test case #800/2803" severity error;
    assert SOL = '0' report "Error in test case #800/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #801/2803" severity error;
    assert SOR = '1' report "Error in test case #801/2803" severity error;
    assert SOL = '0' report "Error in test case #801/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #802/2803" severity error;
    assert SOR = '1' report "Error in test case #802/2803" severity error;
    assert SOL = '0' report "Error in test case #802/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "001";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #803/2803" severity error;
    assert SOR = '1' report "Error in test case #803/2803" severity error;
    assert SOL = '0' report "Error in test case #803/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #804/2803" severity error;
    assert SOR = '1' report "Error in test case #804/2803" severity error;
    assert SOL = '0' report "Error in test case #804/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #805/2803" severity error;
    assert SOR = '1' report "Error in test case #805/2803" severity error;
    assert SOL = '0' report "Error in test case #805/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #806/2803" severity error;
    assert SOR = '1' report "Error in test case #806/2803" severity error;
    assert SOL = '0' report "Error in test case #806/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #807/2803" severity error;
    assert SOR = '1' report "Error in test case #807/2803" severity error;
    assert SOL = '0' report "Error in test case #807/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #808/2803" severity error;
    assert SOR = '0' report "Error in test case #808/2803" severity error;
    assert SOL = '1' report "Error in test case #808/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #809/2803" severity error;
    assert SOR = '0' report "Error in test case #809/2803" severity error;
    assert SOL = '1' report "Error in test case #809/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #810/2803" severity error;
    assert SOR = '0' report "Error in test case #810/2803" severity error;
    assert SOL = '1' report "Error in test case #810/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #811/2803" severity error;
    assert SOR = '0' report "Error in test case #811/2803" severity error;
    assert SOL = '1' report "Error in test case #811/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #812/2803" severity error;
    assert SOR = '0' report "Error in test case #812/2803" severity error;
    assert SOL = '0' report "Error in test case #812/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #813/2803" severity error;
    assert SOR = '0' report "Error in test case #813/2803" severity error;
    assert SOL = '0' report "Error in test case #813/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #814/2803" severity error;
    assert SOR = '0' report "Error in test case #814/2803" severity error;
    assert SOL = '0' report "Error in test case #814/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #815/2803" severity error;
    assert SOR = '0' report "Error in test case #815/2803" severity error;
    assert SOL = '0' report "Error in test case #815/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #816/2803" severity error;
    assert SOR = '1' report "Error in test case #816/2803" severity error;
    assert SOL = '0' report "Error in test case #816/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #817/2803" severity error;
    assert SOR = '1' report "Error in test case #817/2803" severity error;
    assert SOL = '0' report "Error in test case #817/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #818/2803" severity error;
    assert SOR = '1' report "Error in test case #818/2803" severity error;
    assert SOL = '0' report "Error in test case #818/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #819/2803" severity error;
    assert SOR = '1' report "Error in test case #819/2803" severity error;
    assert SOL = '0' report "Error in test case #819/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #820/2803" severity error;
    assert SOR = '1' report "Error in test case #820/2803" severity error;
    assert SOL = '0' report "Error in test case #820/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #821/2803" severity error;
    assert SOR = '1' report "Error in test case #821/2803" severity error;
    assert SOL = '1' report "Error in test case #821/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #822/2803" severity error;
    assert SOR = '1' report "Error in test case #822/2803" severity error;
    assert SOL = '1' report "Error in test case #822/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #823/2803" severity error;
    assert SOR = '1' report "Error in test case #823/2803" severity error;
    assert SOL = '1' report "Error in test case #823/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #824/2803" severity error;
    assert SOR = '0' report "Error in test case #824/2803" severity error;
    assert SOL = '1' report "Error in test case #824/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #825/2803" severity error;
    assert SOR = '0' report "Error in test case #825/2803" severity error;
    assert SOL = '1' report "Error in test case #825/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #826/2803" severity error;
    assert SOR = '0' report "Error in test case #826/2803" severity error;
    assert SOL = '1' report "Error in test case #826/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #827/2803" severity error;
    assert SOR = '0' report "Error in test case #827/2803" severity error;
    assert SOL = '1' report "Error in test case #827/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #828/2803" severity error;
    assert SOR = '0' report "Error in test case #828/2803" severity error;
    assert SOL = '1' report "Error in test case #828/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #829/2803" severity error;
    assert SOR = '0' report "Error in test case #829/2803" severity error;
    assert SOL = '1' report "Error in test case #829/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #830/2803" severity error;
    assert SOR = '0' report "Error in test case #830/2803" severity error;
    assert SOL = '1' report "Error in test case #830/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #831/2803" severity error;
    assert SOR = '1' report "Error in test case #831/2803" severity error;
    assert SOL = '1' report "Error in test case #831/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #832/2803" severity error;
    assert SOR = '0' report "Error in test case #832/2803" severity error;
    assert SOL = '1' report "Error in test case #832/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #833/2803" severity error;
    assert SOR = '0' report "Error in test case #833/2803" severity error;
    assert SOL = '1' report "Error in test case #833/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #834/2803" severity error;
    assert SOR = '0' report "Error in test case #834/2803" severity error;
    assert SOL = '1' report "Error in test case #834/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #835/2803" severity error;
    assert SOR = '0' report "Error in test case #835/2803" severity error;
    assert SOL = '1' report "Error in test case #835/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #836/2803" severity error;
    assert SOR = '0' report "Error in test case #836/2803" severity error;
    assert SOL = '1' report "Error in test case #836/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #837/2803" severity error;
    assert SOR = '0' report "Error in test case #837/2803" severity error;
    assert SOL = '1' report "Error in test case #837/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #838/2803" severity error;
    assert SOR = '0' report "Error in test case #838/2803" severity error;
    assert SOL = '1' report "Error in test case #838/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #839/2803" severity error;
    assert SOR = '0' report "Error in test case #839/2803" severity error;
    assert SOL = '1' report "Error in test case #839/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111100" report "Error in test case #840/2803" severity error;
    assert SOR = '0' report "Error in test case #840/2803" severity error;
    assert SOL = '1' report "Error in test case #840/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111100" report "Error in test case #841/2803" severity error;
    assert SOR = '0' report "Error in test case #841/2803" severity error;
    assert SOL = '1' report "Error in test case #841/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111100" report "Error in test case #842/2803" severity error;
    assert SOR = '0' report "Error in test case #842/2803" severity error;
    assert SOL = '1' report "Error in test case #842/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111100" report "Error in test case #843/2803" severity error;
    assert SOR = '0' report "Error in test case #843/2803" severity error;
    assert SOL = '1' report "Error in test case #843/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111100" report "Error in test case #844/2803" severity error;
    assert SOR = '0' report "Error in test case #844/2803" severity error;
    assert SOL = '1' report "Error in test case #844/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #845/2803" severity error;
    assert SOR = '1' report "Error in test case #845/2803" severity error;
    assert SOL = '1' report "Error in test case #845/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #846/2803" severity error;
    assert SOR = '1' report "Error in test case #846/2803" severity error;
    assert SOL = '1' report "Error in test case #846/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #847/2803" severity error;
    assert SOR = '1' report "Error in test case #847/2803" severity error;
    assert SOL = '1' report "Error in test case #847/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #848/2803" severity error;
    assert SOR = '1' report "Error in test case #848/2803" severity error;
    assert SOL = '1' report "Error in test case #848/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #849/2803" severity error;
    assert SOR = '1' report "Error in test case #849/2803" severity error;
    assert SOL = '1' report "Error in test case #849/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #850/2803" severity error;
    assert SOR = '1' report "Error in test case #850/2803" severity error;
    assert SOL = '1' report "Error in test case #850/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #851/2803" severity error;
    assert SOR = '1' report "Error in test case #851/2803" severity error;
    assert SOL = '1' report "Error in test case #851/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #852/2803" severity error;
    assert SOR = '1' report "Error in test case #852/2803" severity error;
    assert SOL = '1' report "Error in test case #852/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #853/2803" severity error;
    assert SOR = '0' report "Error in test case #853/2803" severity error;
    assert SOL = '0' report "Error in test case #853/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #854/2803" severity error;
    assert SOR = '0' report "Error in test case #854/2803" severity error;
    assert SOL = '0' report "Error in test case #854/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #855/2803" severity error;
    assert SOR = '0' report "Error in test case #855/2803" severity error;
    assert SOL = '0' report "Error in test case #855/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #856/2803" severity error;
    assert SOR = '0' report "Error in test case #856/2803" severity error;
    assert SOL = '0' report "Error in test case #856/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #857/2803" severity error;
    assert SOR = '0' report "Error in test case #857/2803" severity error;
    assert SOL = '0' report "Error in test case #857/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #858/2803" severity error;
    assert SOR = '0' report "Error in test case #858/2803" severity error;
    assert SOL = '0' report "Error in test case #858/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #859/2803" severity error;
    assert SOR = '0' report "Error in test case #859/2803" severity error;
    assert SOL = '0' report "Error in test case #859/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #860/2803" severity error;
    assert SOR = '0' report "Error in test case #860/2803" severity error;
    assert SOL = '0' report "Error in test case #860/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #861/2803" severity error;
    assert SOR = '0' report "Error in test case #861/2803" severity error;
    assert SOL = '0' report "Error in test case #861/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #862/2803" severity error;
    assert SOR = '0' report "Error in test case #862/2803" severity error;
    assert SOL = '0' report "Error in test case #862/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #863/2803" severity error;
    assert SOR = '0' report "Error in test case #863/2803" severity error;
    assert SOL = '0' report "Error in test case #863/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #864/2803" severity error;
    assert SOR = '0' report "Error in test case #864/2803" severity error;
    assert SOL = '0' report "Error in test case #864/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #865/2803" severity error;
    assert SOR = '0' report "Error in test case #865/2803" severity error;
    assert SOL = '0' report "Error in test case #865/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #866/2803" severity error;
    assert SOR = '0' report "Error in test case #866/2803" severity error;
    assert SOL = '0' report "Error in test case #866/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #867/2803" severity error;
    assert SOR = '0' report "Error in test case #867/2803" severity error;
    assert SOL = '0' report "Error in test case #867/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #868/2803" severity error;
    assert SOR = '0' report "Error in test case #868/2803" severity error;
    assert SOL = '0' report "Error in test case #868/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #869/2803" severity error;
    assert SOR = '0' report "Error in test case #869/2803" severity error;
    assert SOL = '0' report "Error in test case #869/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #870/2803" severity error;
    assert SOR = '0' report "Error in test case #870/2803" severity error;
    assert SOL = '0' report "Error in test case #870/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #871/2803" severity error;
    assert SOR = '0' report "Error in test case #871/2803" severity error;
    assert SOL = '0' report "Error in test case #871/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #872/2803" severity error;
    assert SOR = '0' report "Error in test case #872/2803" severity error;
    assert SOL = '0' report "Error in test case #872/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #873/2803" severity error;
    assert SOR = '0' report "Error in test case #873/2803" severity error;
    assert SOL = '0' report "Error in test case #873/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #874/2803" severity error;
    assert SOR = '0' report "Error in test case #874/2803" severity error;
    assert SOL = '0' report "Error in test case #874/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #875/2803" severity error;
    assert SOR = '0' report "Error in test case #875/2803" severity error;
    assert SOL = '0' report "Error in test case #875/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #876/2803" severity error;
    assert SOR = '0' report "Error in test case #876/2803" severity error;
    assert SOL = '0' report "Error in test case #876/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #877/2803" severity error;
    assert SOR = '0' report "Error in test case #877/2803" severity error;
    assert SOL = '0' report "Error in test case #877/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #878/2803" severity error;
    assert SOR = '0' report "Error in test case #878/2803" severity error;
    assert SOL = '0' report "Error in test case #878/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #879/2803" severity error;
    assert SOR = '0' report "Error in test case #879/2803" severity error;
    assert SOL = '0' report "Error in test case #879/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #880/2803" severity error;
    assert SOR = '0' report "Error in test case #880/2803" severity error;
    assert SOL = '0' report "Error in test case #880/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #881/2803" severity error;
    assert SOR = '0' report "Error in test case #881/2803" severity error;
    assert SOL = '0' report "Error in test case #881/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #882/2803" severity error;
    assert SOR = '0' report "Error in test case #882/2803" severity error;
    assert SOL = '0' report "Error in test case #882/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #883/2803" severity error;
    assert SOR = '0' report "Error in test case #883/2803" severity error;
    assert SOL = '0' report "Error in test case #883/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #884/2803" severity error;
    assert SOR = '0' report "Error in test case #884/2803" severity error;
    assert SOL = '0' report "Error in test case #884/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #885/2803" severity error;
    assert SOR = '0' report "Error in test case #885/2803" severity error;
    assert SOL = '0' report "Error in test case #885/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #886/2803" severity error;
    assert SOR = '0' report "Error in test case #886/2803" severity error;
    assert SOL = '0' report "Error in test case #886/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #887/2803" severity error;
    assert SOR = '0' report "Error in test case #887/2803" severity error;
    assert SOL = '0' report "Error in test case #887/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #888/2803" severity error;
    assert SOR = '0' report "Error in test case #888/2803" severity error;
    assert SOL = '0' report "Error in test case #888/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #889/2803" severity error;
    assert SOR = '0' report "Error in test case #889/2803" severity error;
    assert SOL = '0' report "Error in test case #889/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #890/2803" severity error;
    assert SOR = '0' report "Error in test case #890/2803" severity error;
    assert SOL = '0' report "Error in test case #890/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #891/2803" severity error;
    assert SOR = '0' report "Error in test case #891/2803" severity error;
    assert SOL = '0' report "Error in test case #891/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #892/2803" severity error;
    assert SOR = '0' report "Error in test case #892/2803" severity error;
    assert SOL = '0' report "Error in test case #892/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #893/2803" severity error;
    assert SOR = '0' report "Error in test case #893/2803" severity error;
    assert SOL = '0' report "Error in test case #893/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #894/2803" severity error;
    assert SOR = '0' report "Error in test case #894/2803" severity error;
    assert SOL = '0' report "Error in test case #894/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #895/2803" severity error;
    assert SOR = '0' report "Error in test case #895/2803" severity error;
    assert SOL = '0' report "Error in test case #895/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #896/2803" severity error;
    assert SOR = '1' report "Error in test case #896/2803" severity error;
    assert SOL = '1' report "Error in test case #896/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #897/2803" severity error;
    assert SOR = '1' report "Error in test case #897/2803" severity error;
    assert SOL = '1' report "Error in test case #897/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #898/2803" severity error;
    assert SOR = '1' report "Error in test case #898/2803" severity error;
    assert SOL = '1' report "Error in test case #898/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #899/2803" severity error;
    assert SOR = '0' report "Error in test case #899/2803" severity error;
    assert SOL = '0' report "Error in test case #899/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #900/2803" severity error;
    assert SOR = '0' report "Error in test case #900/2803" severity error;
    assert SOL = '0' report "Error in test case #900/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #901/2803" severity error;
    assert SOR = '0' report "Error in test case #901/2803" severity error;
    assert SOL = '0' report "Error in test case #901/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #902/2803" severity error;
    assert SOR = '0' report "Error in test case #902/2803" severity error;
    assert SOL = '0' report "Error in test case #902/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #903/2803" severity error;
    assert SOR = '0' report "Error in test case #903/2803" severity error;
    assert SOL = '0' report "Error in test case #903/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #904/2803" severity error;
    assert SOR = '0' report "Error in test case #904/2803" severity error;
    assert SOL = '0' report "Error in test case #904/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #905/2803" severity error;
    assert SOR = '0' report "Error in test case #905/2803" severity error;
    assert SOL = '0' report "Error in test case #905/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #906/2803" severity error;
    assert SOR = '0' report "Error in test case #906/2803" severity error;
    assert SOL = '0' report "Error in test case #906/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #907/2803" severity error;
    assert SOR = '0' report "Error in test case #907/2803" severity error;
    assert SOL = '0' report "Error in test case #907/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #908/2803" severity error;
    assert SOR = '0' report "Error in test case #908/2803" severity error;
    assert SOL = '0' report "Error in test case #908/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #909/2803" severity error;
    assert SOR = '0' report "Error in test case #909/2803" severity error;
    assert SOL = '0' report "Error in test case #909/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #910/2803" severity error;
    assert SOR = '0' report "Error in test case #910/2803" severity error;
    assert SOL = '0' report "Error in test case #910/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #911/2803" severity error;
    assert SOR = '0' report "Error in test case #911/2803" severity error;
    assert SOL = '0' report "Error in test case #911/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #912/2803" severity error;
    assert SOR = '1' report "Error in test case #912/2803" severity error;
    assert SOL = '0' report "Error in test case #912/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #913/2803" severity error;
    assert SOR = '1' report "Error in test case #913/2803" severity error;
    assert SOL = '0' report "Error in test case #913/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #914/2803" severity error;
    assert SOR = '1' report "Error in test case #914/2803" severity error;
    assert SOL = '0' report "Error in test case #914/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #915/2803" severity error;
    assert SOR = '1' report "Error in test case #915/2803" severity error;
    assert SOL = '0' report "Error in test case #915/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #916/2803" severity error;
    assert SOR = '1' report "Error in test case #916/2803" severity error;
    assert SOL = '0' report "Error in test case #916/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #917/2803" severity error;
    assert SOR = '1' report "Error in test case #917/2803" severity error;
    assert SOL = '0' report "Error in test case #917/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #918/2803" severity error;
    assert SOR = '1' report "Error in test case #918/2803" severity error;
    assert SOL = '0' report "Error in test case #918/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #919/2803" severity error;
    assert SOR = '1' report "Error in test case #919/2803" severity error;
    assert SOL = '0' report "Error in test case #919/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #920/2803" severity error;
    assert SOR = '1' report "Error in test case #920/2803" severity error;
    assert SOL = '0' report "Error in test case #920/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #921/2803" severity error;
    assert SOR = '1' report "Error in test case #921/2803" severity error;
    assert SOL = '0' report "Error in test case #921/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #922/2803" severity error;
    assert SOR = '1' report "Error in test case #922/2803" severity error;
    assert SOL = '0' report "Error in test case #922/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #923/2803" severity error;
    assert SOR = '1' report "Error in test case #923/2803" severity error;
    assert SOL = '0' report "Error in test case #923/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #924/2803" severity error;
    assert SOR = '1' report "Error in test case #924/2803" severity error;
    assert SOL = '0' report "Error in test case #924/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #925/2803" severity error;
    assert SOR = '1' report "Error in test case #925/2803" severity error;
    assert SOL = '0' report "Error in test case #925/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #926/2803" severity error;
    assert SOR = '1' report "Error in test case #926/2803" severity error;
    assert SOL = '0' report "Error in test case #926/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #927/2803" severity error;
    assert SOR = '1' report "Error in test case #927/2803" severity error;
    assert SOL = '0' report "Error in test case #927/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #928/2803" severity error;
    assert SOR = '0' report "Error in test case #928/2803" severity error;
    assert SOL = '0' report "Error in test case #928/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #929/2803" severity error;
    assert SOR = '0' report "Error in test case #929/2803" severity error;
    assert SOL = '0' report "Error in test case #929/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #930/2803" severity error;
    assert SOR = '0' report "Error in test case #930/2803" severity error;
    assert SOL = '0' report "Error in test case #930/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #931/2803" severity error;
    assert SOR = '0' report "Error in test case #931/2803" severity error;
    assert SOL = '0' report "Error in test case #931/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #932/2803" severity error;
    assert SOR = '0' report "Error in test case #932/2803" severity error;
    assert SOL = '0' report "Error in test case #932/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #933/2803" severity error;
    assert SOR = '0' report "Error in test case #933/2803" severity error;
    assert SOL = '0' report "Error in test case #933/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #934/2803" severity error;
    assert SOR = '0' report "Error in test case #934/2803" severity error;
    assert SOL = '0' report "Error in test case #934/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #935/2803" severity error;
    assert SOR = '0' report "Error in test case #935/2803" severity error;
    assert SOL = '0' report "Error in test case #935/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001101" report "Error in test case #936/2803" severity error;
    assert SOR = '1' report "Error in test case #936/2803" severity error;
    assert SOL = '0' report "Error in test case #936/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001101" report "Error in test case #937/2803" severity error;
    assert SOR = '1' report "Error in test case #937/2803" severity error;
    assert SOL = '0' report "Error in test case #937/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001101" report "Error in test case #938/2803" severity error;
    assert SOR = '1' report "Error in test case #938/2803" severity error;
    assert SOL = '0' report "Error in test case #938/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001101" report "Error in test case #939/2803" severity error;
    assert SOR = '1' report "Error in test case #939/2803" severity error;
    assert SOL = '0' report "Error in test case #939/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001101" report "Error in test case #940/2803" severity error;
    assert SOR = '1' report "Error in test case #940/2803" severity error;
    assert SOL = '0' report "Error in test case #940/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001101" report "Error in test case #941/2803" severity error;
    assert SOR = '1' report "Error in test case #941/2803" severity error;
    assert SOL = '0' report "Error in test case #941/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001101" report "Error in test case #942/2803" severity error;
    assert SOR = '1' report "Error in test case #942/2803" severity error;
    assert SOL = '0' report "Error in test case #942/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001101" report "Error in test case #943/2803" severity error;
    assert SOR = '1' report "Error in test case #943/2803" severity error;
    assert SOL = '0' report "Error in test case #943/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011011" report "Error in test case #944/2803" severity error;
    assert SOR = '1' report "Error in test case #944/2803" severity error;
    assert SOL = '0' report "Error in test case #944/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011011" report "Error in test case #945/2803" severity error;
    assert SOR = '1' report "Error in test case #945/2803" severity error;
    assert SOL = '0' report "Error in test case #945/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011011" report "Error in test case #946/2803" severity error;
    assert SOR = '1' report "Error in test case #946/2803" severity error;
    assert SOL = '0' report "Error in test case #946/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011011" report "Error in test case #947/2803" severity error;
    assert SOR = '1' report "Error in test case #947/2803" severity error;
    assert SOL = '0' report "Error in test case #947/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011011" report "Error in test case #948/2803" severity error;
    assert SOR = '1' report "Error in test case #948/2803" severity error;
    assert SOL = '0' report "Error in test case #948/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011011" report "Error in test case #949/2803" severity error;
    assert SOR = '1' report "Error in test case #949/2803" severity error;
    assert SOL = '0' report "Error in test case #949/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011011" report "Error in test case #950/2803" severity error;
    assert SOR = '1' report "Error in test case #950/2803" severity error;
    assert SOL = '0' report "Error in test case #950/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011011" report "Error in test case #951/2803" severity error;
    assert SOR = '1' report "Error in test case #951/2803" severity error;
    assert SOL = '0' report "Error in test case #951/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00110111" report "Error in test case #952/2803" severity error;
    assert SOR = '1' report "Error in test case #952/2803" severity error;
    assert SOL = '0' report "Error in test case #952/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00110111" report "Error in test case #953/2803" severity error;
    assert SOR = '1' report "Error in test case #953/2803" severity error;
    assert SOL = '0' report "Error in test case #953/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00110111" report "Error in test case #954/2803" severity error;
    assert SOR = '1' report "Error in test case #954/2803" severity error;
    assert SOL = '0' report "Error in test case #954/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00110111" report "Error in test case #955/2803" severity error;
    assert SOR = '1' report "Error in test case #955/2803" severity error;
    assert SOL = '0' report "Error in test case #955/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00110111" report "Error in test case #956/2803" severity error;
    assert SOR = '1' report "Error in test case #956/2803" severity error;
    assert SOL = '0' report "Error in test case #956/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00110111" report "Error in test case #957/2803" severity error;
    assert SOR = '1' report "Error in test case #957/2803" severity error;
    assert SOL = '0' report "Error in test case #957/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00110111" report "Error in test case #958/2803" severity error;
    assert SOR = '1' report "Error in test case #958/2803" severity error;
    assert SOL = '0' report "Error in test case #958/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00110111" report "Error in test case #959/2803" severity error;
    assert SOR = '1' report "Error in test case #959/2803" severity error;
    assert SOL = '0' report "Error in test case #959/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01101110" report "Error in test case #960/2803" severity error;
    assert SOR = '0' report "Error in test case #960/2803" severity error;
    assert SOL = '0' report "Error in test case #960/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01101110" report "Error in test case #961/2803" severity error;
    assert SOR = '0' report "Error in test case #961/2803" severity error;
    assert SOL = '0' report "Error in test case #961/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01101110" report "Error in test case #962/2803" severity error;
    assert SOR = '0' report "Error in test case #962/2803" severity error;
    assert SOL = '0' report "Error in test case #962/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01101110" report "Error in test case #963/2803" severity error;
    assert SOR = '0' report "Error in test case #963/2803" severity error;
    assert SOL = '0' report "Error in test case #963/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01101110" report "Error in test case #964/2803" severity error;
    assert SOR = '0' report "Error in test case #964/2803" severity error;
    assert SOL = '0' report "Error in test case #964/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #965/2803" severity error;
    assert SOR = '1' report "Error in test case #965/2803" severity error;
    assert SOL = '1' report "Error in test case #965/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #966/2803" severity error;
    assert SOR = '1' report "Error in test case #966/2803" severity error;
    assert SOL = '1' report "Error in test case #966/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #967/2803" severity error;
    assert SOR = '1' report "Error in test case #967/2803" severity error;
    assert SOL = '1' report "Error in test case #967/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #968/2803" severity error;
    assert SOR = '1' report "Error in test case #968/2803" severity error;
    assert SOL = '1' report "Error in test case #968/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #969/2803" severity error;
    assert SOR = '1' report "Error in test case #969/2803" severity error;
    assert SOL = '1' report "Error in test case #969/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #970/2803" severity error;
    assert SOR = '1' report "Error in test case #970/2803" severity error;
    assert SOL = '1' report "Error in test case #970/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #971/2803" severity error;
    assert SOR = '1' report "Error in test case #971/2803" severity error;
    assert SOL = '1' report "Error in test case #971/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #972/2803" severity error;
    assert SOR = '1' report "Error in test case #972/2803" severity error;
    assert SOL = '1' report "Error in test case #972/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #973/2803" severity error;
    assert SOR = '1' report "Error in test case #973/2803" severity error;
    assert SOL = '1' report "Error in test case #973/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #974/2803" severity error;
    assert SOR = '1' report "Error in test case #974/2803" severity error;
    assert SOL = '1' report "Error in test case #974/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #975/2803" severity error;
    assert SOR = '1' report "Error in test case #975/2803" severity error;
    assert SOL = '1' report "Error in test case #975/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #976/2803" severity error;
    assert SOR = '1' report "Error in test case #976/2803" severity error;
    assert SOL = '1' report "Error in test case #976/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #977/2803" severity error;
    assert SOR = '1' report "Error in test case #977/2803" severity error;
    assert SOL = '1' report "Error in test case #977/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #978/2803" severity error;
    assert SOR = '1' report "Error in test case #978/2803" severity error;
    assert SOL = '1' report "Error in test case #978/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #979/2803" severity error;
    assert SOR = '1' report "Error in test case #979/2803" severity error;
    assert SOL = '1' report "Error in test case #979/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #980/2803" severity error;
    assert SOR = '1' report "Error in test case #980/2803" severity error;
    assert SOL = '1' report "Error in test case #980/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #981/2803" severity error;
    assert SOR = '1' report "Error in test case #981/2803" severity error;
    assert SOL = '1' report "Error in test case #981/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #982/2803" severity error;
    assert SOR = '1' report "Error in test case #982/2803" severity error;
    assert SOL = '1' report "Error in test case #982/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #983/2803" severity error;
    assert SOR = '1' report "Error in test case #983/2803" severity error;
    assert SOL = '1' report "Error in test case #983/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #984/2803" severity error;
    assert SOR = '0' report "Error in test case #984/2803" severity error;
    assert SOL = '1' report "Error in test case #984/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #985/2803" severity error;
    assert SOR = '0' report "Error in test case #985/2803" severity error;
    assert SOL = '1' report "Error in test case #985/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #986/2803" severity error;
    assert SOR = '0' report "Error in test case #986/2803" severity error;
    assert SOL = '1' report "Error in test case #986/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #987/2803" severity error;
    assert SOR = '0' report "Error in test case #987/2803" severity error;
    assert SOL = '1' report "Error in test case #987/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #988/2803" severity error;
    assert SOR = '0' report "Error in test case #988/2803" severity error;
    assert SOL = '1' report "Error in test case #988/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #989/2803" severity error;
    assert SOR = '0' report "Error in test case #989/2803" severity error;
    assert SOL = '1' report "Error in test case #989/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #990/2803" severity error;
    assert SOR = '0' report "Error in test case #990/2803" severity error;
    assert SOL = '1' report "Error in test case #990/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #991/2803" severity error;
    assert SOR = '0' report "Error in test case #991/2803" severity error;
    assert SOL = '1' report "Error in test case #991/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #992/2803" severity error;
    assert SOR = '1' report "Error in test case #992/2803" severity error;
    assert SOL = '1' report "Error in test case #992/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #993/2803" severity error;
    assert SOR = '1' report "Error in test case #993/2803" severity error;
    assert SOL = '1' report "Error in test case #993/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #994/2803" severity error;
    assert SOR = '1' report "Error in test case #994/2803" severity error;
    assert SOL = '1' report "Error in test case #994/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #995/2803" severity error;
    assert SOR = '1' report "Error in test case #995/2803" severity error;
    assert SOL = '1' report "Error in test case #995/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #996/2803" severity error;
    assert SOR = '1' report "Error in test case #996/2803" severity error;
    assert SOL = '1' report "Error in test case #996/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #997/2803" severity error;
    assert SOR = '1' report "Error in test case #997/2803" severity error;
    assert SOL = '1' report "Error in test case #997/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #998/2803" severity error;
    assert SOR = '1' report "Error in test case #998/2803" severity error;
    assert SOL = '1' report "Error in test case #998/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #999/2803" severity error;
    assert SOR = '1' report "Error in test case #999/2803" severity error;
    assert SOL = '1' report "Error in test case #999/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1000/2803" severity error;
    assert SOR = '1' report "Error in test case #1000/2803" severity error;
    assert SOL = '1' report "Error in test case #1000/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1001/2803" severity error;
    assert SOR = '1' report "Error in test case #1001/2803" severity error;
    assert SOL = '1' report "Error in test case #1001/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1002/2803" severity error;
    assert SOR = '1' report "Error in test case #1002/2803" severity error;
    assert SOL = '1' report "Error in test case #1002/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1003/2803" severity error;
    assert SOR = '1' report "Error in test case #1003/2803" severity error;
    assert SOL = '1' report "Error in test case #1003/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1004/2803" severity error;
    assert SOR = '1' report "Error in test case #1004/2803" severity error;
    assert SOL = '1' report "Error in test case #1004/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1005/2803" severity error;
    assert SOR = '1' report "Error in test case #1005/2803" severity error;
    assert SOL = '1' report "Error in test case #1005/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1006/2803" severity error;
    assert SOR = '1' report "Error in test case #1006/2803" severity error;
    assert SOL = '1' report "Error in test case #1006/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1007/2803" severity error;
    assert SOR = '1' report "Error in test case #1007/2803" severity error;
    assert SOL = '1' report "Error in test case #1007/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1008/2803" severity error;
    assert SOR = '1' report "Error in test case #1008/2803" severity error;
    assert SOL = '1' report "Error in test case #1008/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1009/2803" severity error;
    assert SOR = '1' report "Error in test case #1009/2803" severity error;
    assert SOL = '1' report "Error in test case #1009/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1010/2803" severity error;
    assert SOR = '1' report "Error in test case #1010/2803" severity error;
    assert SOL = '1' report "Error in test case #1010/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1011/2803" severity error;
    assert SOR = '1' report "Error in test case #1011/2803" severity error;
    assert SOL = '1' report "Error in test case #1011/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1012/2803" severity error;
    assert SOR = '0' report "Error in test case #1012/2803" severity error;
    assert SOL = '0' report "Error in test case #1012/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1013/2803" severity error;
    assert SOR = '0' report "Error in test case #1013/2803" severity error;
    assert SOL = '0' report "Error in test case #1013/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1014/2803" severity error;
    assert SOR = '0' report "Error in test case #1014/2803" severity error;
    assert SOL = '0' report "Error in test case #1014/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1015/2803" severity error;
    assert SOR = '0' report "Error in test case #1015/2803" severity error;
    assert SOL = '0' report "Error in test case #1015/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1016/2803" severity error;
    assert SOR = '1' report "Error in test case #1016/2803" severity error;
    assert SOL = '0' report "Error in test case #1016/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1017/2803" severity error;
    assert SOR = '1' report "Error in test case #1017/2803" severity error;
    assert SOL = '0' report "Error in test case #1017/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1018/2803" severity error;
    assert SOR = '1' report "Error in test case #1018/2803" severity error;
    assert SOL = '0' report "Error in test case #1018/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1019/2803" severity error;
    assert SOR = '1' report "Error in test case #1019/2803" severity error;
    assert SOL = '0' report "Error in test case #1019/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1020/2803" severity error;
    assert SOR = '1' report "Error in test case #1020/2803" severity error;
    assert SOL = '0' report "Error in test case #1020/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1021/2803" severity error;
    assert SOR = '1' report "Error in test case #1021/2803" severity error;
    assert SOL = '0' report "Error in test case #1021/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1022/2803" severity error;
    assert SOR = '1' report "Error in test case #1022/2803" severity error;
    assert SOL = '0' report "Error in test case #1022/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1023/2803" severity error;
    assert SOR = '1' report "Error in test case #1023/2803" severity error;
    assert SOL = '0' report "Error in test case #1023/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1024/2803" severity error;
    assert SOR = '1' report "Error in test case #1024/2803" severity error;
    assert SOL = '0' report "Error in test case #1024/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1025/2803" severity error;
    assert SOR = '1' report "Error in test case #1025/2803" severity error;
    assert SOL = '0' report "Error in test case #1025/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1026/2803" severity error;
    assert SOR = '1' report "Error in test case #1026/2803" severity error;
    assert SOL = '0' report "Error in test case #1026/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1027/2803" severity error;
    assert SOR = '1' report "Error in test case #1027/2803" severity error;
    assert SOL = '0' report "Error in test case #1027/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1028/2803" severity error;
    assert SOR = '1' report "Error in test case #1028/2803" severity error;
    assert SOL = '0' report "Error in test case #1028/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1029/2803" severity error;
    assert SOR = '1' report "Error in test case #1029/2803" severity error;
    assert SOL = '0' report "Error in test case #1029/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1030/2803" severity error;
    assert SOR = '1' report "Error in test case #1030/2803" severity error;
    assert SOL = '0' report "Error in test case #1030/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1031/2803" severity error;
    assert SOR = '1' report "Error in test case #1031/2803" severity error;
    assert SOL = '0' report "Error in test case #1031/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1032/2803" severity error;
    assert SOR = '1' report "Error in test case #1032/2803" severity error;
    assert SOL = '0' report "Error in test case #1032/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1033/2803" severity error;
    assert SOR = '1' report "Error in test case #1033/2803" severity error;
    assert SOL = '0' report "Error in test case #1033/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1034/2803" severity error;
    assert SOR = '1' report "Error in test case #1034/2803" severity error;
    assert SOL = '0' report "Error in test case #1034/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1035/2803" severity error;
    assert SOR = '1' report "Error in test case #1035/2803" severity error;
    assert SOL = '0' report "Error in test case #1035/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1036/2803" severity error;
    assert SOR = '1' report "Error in test case #1036/2803" severity error;
    assert SOL = '0' report "Error in test case #1036/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1037/2803" severity error;
    assert SOR = '1' report "Error in test case #1037/2803" severity error;
    assert SOL = '0' report "Error in test case #1037/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1038/2803" severity error;
    assert SOR = '1' report "Error in test case #1038/2803" severity error;
    assert SOL = '0' report "Error in test case #1038/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1039/2803" severity error;
    assert SOR = '1' report "Error in test case #1039/2803" severity error;
    assert SOL = '0' report "Error in test case #1039/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #1040/2803" severity error;
    assert SOR = '1' report "Error in test case #1040/2803" severity error;
    assert SOL = '0' report "Error in test case #1040/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #1041/2803" severity error;
    assert SOR = '1' report "Error in test case #1041/2803" severity error;
    assert SOL = '0' report "Error in test case #1041/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #1042/2803" severity error;
    assert SOR = '1' report "Error in test case #1042/2803" severity error;
    assert SOL = '0' report "Error in test case #1042/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #1043/2803" severity error;
    assert SOR = '1' report "Error in test case #1043/2803" severity error;
    assert SOL = '0' report "Error in test case #1043/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #1044/2803" severity error;
    assert SOR = '1' report "Error in test case #1044/2803" severity error;
    assert SOL = '0' report "Error in test case #1044/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #1045/2803" severity error;
    assert SOR = '1' report "Error in test case #1045/2803" severity error;
    assert SOL = '0' report "Error in test case #1045/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #1046/2803" severity error;
    assert SOR = '1' report "Error in test case #1046/2803" severity error;
    assert SOL = '0' report "Error in test case #1046/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001111" report "Error in test case #1047/2803" severity error;
    assert SOR = '1' report "Error in test case #1047/2803" severity error;
    assert SOL = '0' report "Error in test case #1047/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #1048/2803" severity error;
    assert SOR = '1' report "Error in test case #1048/2803" severity error;
    assert SOL = '0' report "Error in test case #1048/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #1049/2803" severity error;
    assert SOR = '1' report "Error in test case #1049/2803" severity error;
    assert SOL = '0' report "Error in test case #1049/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #1050/2803" severity error;
    assert SOR = '1' report "Error in test case #1050/2803" severity error;
    assert SOL = '0' report "Error in test case #1050/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #1051/2803" severity error;
    assert SOR = '1' report "Error in test case #1051/2803" severity error;
    assert SOL = '0' report "Error in test case #1051/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #1052/2803" severity error;
    assert SOR = '1' report "Error in test case #1052/2803" severity error;
    assert SOL = '0' report "Error in test case #1052/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #1053/2803" severity error;
    assert SOR = '1' report "Error in test case #1053/2803" severity error;
    assert SOL = '0' report "Error in test case #1053/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #1054/2803" severity error;
    assert SOR = '1' report "Error in test case #1054/2803" severity error;
    assert SOL = '0' report "Error in test case #1054/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00011111" report "Error in test case #1055/2803" severity error;
    assert SOR = '1' report "Error in test case #1055/2803" severity error;
    assert SOL = '0' report "Error in test case #1055/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #1056/2803" severity error;
    assert SOR = '1' report "Error in test case #1056/2803" severity error;
    assert SOL = '0' report "Error in test case #1056/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #1057/2803" severity error;
    assert SOR = '1' report "Error in test case #1057/2803" severity error;
    assert SOL = '0' report "Error in test case #1057/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #1058/2803" severity error;
    assert SOR = '1' report "Error in test case #1058/2803" severity error;
    assert SOL = '0' report "Error in test case #1058/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #1059/2803" severity error;
    assert SOR = '1' report "Error in test case #1059/2803" severity error;
    assert SOL = '0' report "Error in test case #1059/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #1060/2803" severity error;
    assert SOR = '1' report "Error in test case #1060/2803" severity error;
    assert SOL = '0' report "Error in test case #1060/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #1061/2803" severity error;
    assert SOR = '1' report "Error in test case #1061/2803" severity error;
    assert SOL = '0' report "Error in test case #1061/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #1062/2803" severity error;
    assert SOR = '1' report "Error in test case #1062/2803" severity error;
    assert SOL = '0' report "Error in test case #1062/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00111111" report "Error in test case #1063/2803" severity error;
    assert SOR = '1' report "Error in test case #1063/2803" severity error;
    assert SOL = '0' report "Error in test case #1063/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #1064/2803" severity error;
    assert SOR = '1' report "Error in test case #1064/2803" severity error;
    assert SOL = '0' report "Error in test case #1064/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #1065/2803" severity error;
    assert SOR = '1' report "Error in test case #1065/2803" severity error;
    assert SOL = '0' report "Error in test case #1065/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #1066/2803" severity error;
    assert SOR = '1' report "Error in test case #1066/2803" severity error;
    assert SOL = '0' report "Error in test case #1066/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #1067/2803" severity error;
    assert SOR = '1' report "Error in test case #1067/2803" severity error;
    assert SOL = '0' report "Error in test case #1067/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #1068/2803" severity error;
    assert SOR = '1' report "Error in test case #1068/2803" severity error;
    assert SOL = '0' report "Error in test case #1068/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #1069/2803" severity error;
    assert SOR = '1' report "Error in test case #1069/2803" severity error;
    assert SOL = '0' report "Error in test case #1069/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #1070/2803" severity error;
    assert SOR = '1' report "Error in test case #1070/2803" severity error;
    assert SOL = '0' report "Error in test case #1070/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "01111111" report "Error in test case #1071/2803" severity error;
    assert SOR = '1' report "Error in test case #1071/2803" severity error;
    assert SOL = '0' report "Error in test case #1071/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1072/2803" severity error;
    assert SOR = '0' report "Error in test case #1072/2803" severity error;
    assert SOL = '1' report "Error in test case #1072/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1073/2803" severity error;
    assert SOR = '0' report "Error in test case #1073/2803" severity error;
    assert SOL = '1' report "Error in test case #1073/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1074/2803" severity error;
    assert SOR = '0' report "Error in test case #1074/2803" severity error;
    assert SOL = '1' report "Error in test case #1074/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1075/2803" severity error;
    assert SOR = '0' report "Error in test case #1075/2803" severity error;
    assert SOL = '1' report "Error in test case #1075/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1076/2803" severity error;
    assert SOR = '0' report "Error in test case #1076/2803" severity error;
    assert SOL = '1' report "Error in test case #1076/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1077/2803" severity error;
    assert SOR = '0' report "Error in test case #1077/2803" severity error;
    assert SOL = '1' report "Error in test case #1077/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1078/2803" severity error;
    assert SOR = '0' report "Error in test case #1078/2803" severity error;
    assert SOL = '1' report "Error in test case #1078/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1079/2803" severity error;
    assert SOR = '0' report "Error in test case #1079/2803" severity error;
    assert SOL = '1' report "Error in test case #1079/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #1080/2803" severity error;
    assert SOR = '1' report "Error in test case #1080/2803" severity error;
    assert SOL = '1' report "Error in test case #1080/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #1081/2803" severity error;
    assert SOR = '1' report "Error in test case #1081/2803" severity error;
    assert SOL = '1' report "Error in test case #1081/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #1082/2803" severity error;
    assert SOR = '1' report "Error in test case #1082/2803" severity error;
    assert SOL = '1' report "Error in test case #1082/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #1083/2803" severity error;
    assert SOR = '1' report "Error in test case #1083/2803" severity error;
    assert SOL = '1' report "Error in test case #1083/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #1084/2803" severity error;
    assert SOR = '1' report "Error in test case #1084/2803" severity error;
    assert SOL = '1' report "Error in test case #1084/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #1085/2803" severity error;
    assert SOR = '1' report "Error in test case #1085/2803" severity error;
    assert SOL = '1' report "Error in test case #1085/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111101" report "Error in test case #1086/2803" severity error;
    assert SOR = '1' report "Error in test case #1086/2803" severity error;
    assert SOL = '1' report "Error in test case #1086/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1087/2803" severity error;
    assert SOR = '0' report "Error in test case #1087/2803" severity error;
    assert SOL = '0' report "Error in test case #1087/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1088/2803" severity error;
    assert SOR = '0' report "Error in test case #1088/2803" severity error;
    assert SOL = '0' report "Error in test case #1088/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1089/2803" severity error;
    assert SOR = '0' report "Error in test case #1089/2803" severity error;
    assert SOL = '0' report "Error in test case #1089/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1090/2803" severity error;
    assert SOR = '0' report "Error in test case #1090/2803" severity error;
    assert SOL = '0' report "Error in test case #1090/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1091/2803" severity error;
    assert SOR = '0' report "Error in test case #1091/2803" severity error;
    assert SOL = '0' report "Error in test case #1091/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1092/2803" severity error;
    assert SOR = '0' report "Error in test case #1092/2803" severity error;
    assert SOL = '0' report "Error in test case #1092/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1093/2803" severity error;
    assert SOR = '0' report "Error in test case #1093/2803" severity error;
    assert SOL = '0' report "Error in test case #1093/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1094/2803" severity error;
    assert SOR = '0' report "Error in test case #1094/2803" severity error;
    assert SOL = '0' report "Error in test case #1094/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1095/2803" severity error;
    assert SOR = '0' report "Error in test case #1095/2803" severity error;
    assert SOL = '0' report "Error in test case #1095/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1096/2803" severity error;
    assert SOR = '0' report "Error in test case #1096/2803" severity error;
    assert SOL = '0' report "Error in test case #1096/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1097/2803" severity error;
    assert SOR = '0' report "Error in test case #1097/2803" severity error;
    assert SOL = '0' report "Error in test case #1097/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1098/2803" severity error;
    assert SOR = '0' report "Error in test case #1098/2803" severity error;
    assert SOL = '0' report "Error in test case #1098/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1099/2803" severity error;
    assert SOR = '0' report "Error in test case #1099/2803" severity error;
    assert SOL = '0' report "Error in test case #1099/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1100/2803" severity error;
    assert SOR = '0' report "Error in test case #1100/2803" severity error;
    assert SOL = '0' report "Error in test case #1100/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1101/2803" severity error;
    assert SOR = '0' report "Error in test case #1101/2803" severity error;
    assert SOL = '0' report "Error in test case #1101/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1102/2803" severity error;
    assert SOR = '0' report "Error in test case #1102/2803" severity error;
    assert SOL = '0' report "Error in test case #1102/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1103/2803" severity error;
    assert SOR = '0' report "Error in test case #1103/2803" severity error;
    assert SOL = '0' report "Error in test case #1103/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1104/2803" severity error;
    assert SOR = '0' report "Error in test case #1104/2803" severity error;
    assert SOL = '0' report "Error in test case #1104/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1105/2803" severity error;
    assert SOR = '0' report "Error in test case #1105/2803" severity error;
    assert SOL = '0' report "Error in test case #1105/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1106/2803" severity error;
    assert SOR = '0' report "Error in test case #1106/2803" severity error;
    assert SOL = '0' report "Error in test case #1106/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1107/2803" severity error;
    assert SOR = '0' report "Error in test case #1107/2803" severity error;
    assert SOL = '0' report "Error in test case #1107/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1108/2803" severity error;
    assert SOR = '0' report "Error in test case #1108/2803" severity error;
    assert SOL = '0' report "Error in test case #1108/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1109/2803" severity error;
    assert SOR = '0' report "Error in test case #1109/2803" severity error;
    assert SOL = '0' report "Error in test case #1109/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1110/2803" severity error;
    assert SOR = '0' report "Error in test case #1110/2803" severity error;
    assert SOL = '0' report "Error in test case #1110/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1111/2803" severity error;
    assert SOR = '0' report "Error in test case #1111/2803" severity error;
    assert SOL = '0' report "Error in test case #1111/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1112/2803" severity error;
    assert SOR = '1' report "Error in test case #1112/2803" severity error;
    assert SOL = '0' report "Error in test case #1112/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1113/2803" severity error;
    assert SOR = '1' report "Error in test case #1113/2803" severity error;
    assert SOL = '0' report "Error in test case #1113/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1114/2803" severity error;
    assert SOR = '1' report "Error in test case #1114/2803" severity error;
    assert SOL = '0' report "Error in test case #1114/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1115/2803" severity error;
    assert SOR = '1' report "Error in test case #1115/2803" severity error;
    assert SOL = '0' report "Error in test case #1115/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1116/2803" severity error;
    assert SOR = '1' report "Error in test case #1116/2803" severity error;
    assert SOL = '0' report "Error in test case #1116/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1117/2803" severity error;
    assert SOR = '1' report "Error in test case #1117/2803" severity error;
    assert SOL = '0' report "Error in test case #1117/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1118/2803" severity error;
    assert SOR = '1' report "Error in test case #1118/2803" severity error;
    assert SOL = '0' report "Error in test case #1118/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1119/2803" severity error;
    assert SOR = '1' report "Error in test case #1119/2803" severity error;
    assert SOL = '0' report "Error in test case #1119/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1120/2803" severity error;
    assert SOR = '0' report "Error in test case #1120/2803" severity error;
    assert SOL = '0' report "Error in test case #1120/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1121/2803" severity error;
    assert SOR = '0' report "Error in test case #1121/2803" severity error;
    assert SOL = '0' report "Error in test case #1121/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1122/2803" severity error;
    assert SOR = '0' report "Error in test case #1122/2803" severity error;
    assert SOL = '0' report "Error in test case #1122/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1123/2803" severity error;
    assert SOR = '0' report "Error in test case #1123/2803" severity error;
    assert SOL = '0' report "Error in test case #1123/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1124/2803" severity error;
    assert SOR = '0' report "Error in test case #1124/2803" severity error;
    assert SOL = '0' report "Error in test case #1124/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1125/2803" severity error;
    assert SOR = '0' report "Error in test case #1125/2803" severity error;
    assert SOL = '0' report "Error in test case #1125/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1126/2803" severity error;
    assert SOR = '0' report "Error in test case #1126/2803" severity error;
    assert SOL = '0' report "Error in test case #1126/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1127/2803" severity error;
    assert SOR = '0' report "Error in test case #1127/2803" severity error;
    assert SOL = '0' report "Error in test case #1127/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1128/2803" severity error;
    assert SOR = '1' report "Error in test case #1128/2803" severity error;
    assert SOL = '0' report "Error in test case #1128/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1129/2803" severity error;
    assert SOR = '1' report "Error in test case #1129/2803" severity error;
    assert SOL = '0' report "Error in test case #1129/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1130/2803" severity error;
    assert SOR = '1' report "Error in test case #1130/2803" severity error;
    assert SOL = '0' report "Error in test case #1130/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1131/2803" severity error;
    assert SOR = '1' report "Error in test case #1131/2803" severity error;
    assert SOL = '0' report "Error in test case #1131/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1132/2803" severity error;
    assert SOR = '1' report "Error in test case #1132/2803" severity error;
    assert SOL = '0' report "Error in test case #1132/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1133/2803" severity error;
    assert SOR = '1' report "Error in test case #1133/2803" severity error;
    assert SOL = '0' report "Error in test case #1133/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1134/2803" severity error;
    assert SOR = '1' report "Error in test case #1134/2803" severity error;
    assert SOL = '0' report "Error in test case #1134/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1135/2803" severity error;
    assert SOR = '1' report "Error in test case #1135/2803" severity error;
    assert SOL = '0' report "Error in test case #1135/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001011" report "Error in test case #1136/2803" severity error;
    assert SOR = '1' report "Error in test case #1136/2803" severity error;
    assert SOL = '0' report "Error in test case #1136/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001011" report "Error in test case #1137/2803" severity error;
    assert SOR = '1' report "Error in test case #1137/2803" severity error;
    assert SOL = '0' report "Error in test case #1137/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001011" report "Error in test case #1138/2803" severity error;
    assert SOR = '1' report "Error in test case #1138/2803" severity error;
    assert SOL = '0' report "Error in test case #1138/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001011" report "Error in test case #1139/2803" severity error;
    assert SOR = '1' report "Error in test case #1139/2803" severity error;
    assert SOL = '0' report "Error in test case #1139/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00001011" report "Error in test case #1140/2803" severity error;
    assert SOR = '1' report "Error in test case #1140/2803" severity error;
    assert SOL = '0' report "Error in test case #1140/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00001011" report "Error in test case #1141/2803" severity error;
    assert SOR = '1' report "Error in test case #1141/2803" severity error;
    assert SOL = '0' report "Error in test case #1141/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00001011" report "Error in test case #1142/2803" severity error;
    assert SOR = '1' report "Error in test case #1142/2803" severity error;
    assert SOL = '0' report "Error in test case #1142/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00001011" report "Error in test case #1143/2803" severity error;
    assert SOR = '1' report "Error in test case #1143/2803" severity error;
    assert SOL = '0' report "Error in test case #1143/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00010110" report "Error in test case #1144/2803" severity error;
    assert SOR = '0' report "Error in test case #1144/2803" severity error;
    assert SOL = '0' report "Error in test case #1144/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00010110" report "Error in test case #1145/2803" severity error;
    assert SOR = '0' report "Error in test case #1145/2803" severity error;
    assert SOL = '0' report "Error in test case #1145/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00010110" report "Error in test case #1146/2803" severity error;
    assert SOR = '0' report "Error in test case #1146/2803" severity error;
    assert SOL = '0' report "Error in test case #1146/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00010110" report "Error in test case #1147/2803" severity error;
    assert SOR = '0' report "Error in test case #1147/2803" severity error;
    assert SOL = '0' report "Error in test case #1147/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1148/2803" severity error;
    assert SOR = '0' report "Error in test case #1148/2803" severity error;
    assert SOL = '0' report "Error in test case #1148/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1149/2803" severity error;
    assert SOR = '0' report "Error in test case #1149/2803" severity error;
    assert SOL = '0' report "Error in test case #1149/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1150/2803" severity error;
    assert SOR = '0' report "Error in test case #1150/2803" severity error;
    assert SOL = '0' report "Error in test case #1150/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1151/2803" severity error;
    assert SOR = '0' report "Error in test case #1151/2803" severity error;
    assert SOL = '0' report "Error in test case #1151/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1152/2803" severity error;
    assert SOR = '0' report "Error in test case #1152/2803" severity error;
    assert SOL = '0' report "Error in test case #1152/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1153/2803" severity error;
    assert SOR = '0' report "Error in test case #1153/2803" severity error;
    assert SOL = '0' report "Error in test case #1153/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1154/2803" severity error;
    assert SOR = '0' report "Error in test case #1154/2803" severity error;
    assert SOL = '0' report "Error in test case #1154/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1155/2803" severity error;
    assert SOR = '0' report "Error in test case #1155/2803" severity error;
    assert SOL = '0' report "Error in test case #1155/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1156/2803" severity error;
    assert SOR = '0' report "Error in test case #1156/2803" severity error;
    assert SOL = '0' report "Error in test case #1156/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1157/2803" severity error;
    assert SOR = '0' report "Error in test case #1157/2803" severity error;
    assert SOL = '0' report "Error in test case #1157/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1158/2803" severity error;
    assert SOR = '0' report "Error in test case #1158/2803" severity error;
    assert SOL = '0' report "Error in test case #1158/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1159/2803" severity error;
    assert SOR = '0' report "Error in test case #1159/2803" severity error;
    assert SOL = '0' report "Error in test case #1159/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1160/2803" severity error;
    assert SOR = '0' report "Error in test case #1160/2803" severity error;
    assert SOL = '0' report "Error in test case #1160/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1161/2803" severity error;
    assert SOR = '0' report "Error in test case #1161/2803" severity error;
    assert SOL = '0' report "Error in test case #1161/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1162/2803" severity error;
    assert SOR = '0' report "Error in test case #1162/2803" severity error;
    assert SOL = '0' report "Error in test case #1162/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1163/2803" severity error;
    assert SOR = '0' report "Error in test case #1163/2803" severity error;
    assert SOL = '0' report "Error in test case #1163/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1164/2803" severity error;
    assert SOR = '0' report "Error in test case #1164/2803" severity error;
    assert SOL = '0' report "Error in test case #1164/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1165/2803" severity error;
    assert SOR = '0' report "Error in test case #1165/2803" severity error;
    assert SOL = '0' report "Error in test case #1165/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1166/2803" severity error;
    assert SOR = '0' report "Error in test case #1166/2803" severity error;
    assert SOL = '0' report "Error in test case #1166/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1167/2803" severity error;
    assert SOR = '0' report "Error in test case #1167/2803" severity error;
    assert SOL = '0' report "Error in test case #1167/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1168/2803" severity error;
    assert SOR = '1' report "Error in test case #1168/2803" severity error;
    assert SOL = '1' report "Error in test case #1168/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1169/2803" severity error;
    assert SOR = '1' report "Error in test case #1169/2803" severity error;
    assert SOL = '1' report "Error in test case #1169/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1170/2803" severity error;
    assert SOR = '1' report "Error in test case #1170/2803" severity error;
    assert SOL = '1' report "Error in test case #1170/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1171/2803" severity error;
    assert SOR = '1' report "Error in test case #1171/2803" severity error;
    assert SOL = '1' report "Error in test case #1171/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1172/2803" severity error;
    assert SOR = '1' report "Error in test case #1172/2803" severity error;
    assert SOL = '1' report "Error in test case #1172/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1173/2803" severity error;
    assert SOR = '1' report "Error in test case #1173/2803" severity error;
    assert SOL = '1' report "Error in test case #1173/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1174/2803" severity error;
    assert SOR = '1' report "Error in test case #1174/2803" severity error;
    assert SOL = '1' report "Error in test case #1174/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1175/2803" severity error;
    assert SOR = '1' report "Error in test case #1175/2803" severity error;
    assert SOL = '1' report "Error in test case #1175/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1176/2803" severity error;
    assert SOR = '0' report "Error in test case #1176/2803" severity error;
    assert SOL = '1' report "Error in test case #1176/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1177/2803" severity error;
    assert SOR = '0' report "Error in test case #1177/2803" severity error;
    assert SOL = '1' report "Error in test case #1177/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1178/2803" severity error;
    assert SOR = '0' report "Error in test case #1178/2803" severity error;
    assert SOL = '1' report "Error in test case #1178/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1179/2803" severity error;
    assert SOR = '0' report "Error in test case #1179/2803" severity error;
    assert SOL = '1' report "Error in test case #1179/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1180/2803" severity error;
    assert SOR = '0' report "Error in test case #1180/2803" severity error;
    assert SOL = '1' report "Error in test case #1180/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1181/2803" severity error;
    assert SOR = '0' report "Error in test case #1181/2803" severity error;
    assert SOL = '1' report "Error in test case #1181/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111110" report "Error in test case #1182/2803" severity error;
    assert SOR = '0' report "Error in test case #1182/2803" severity error;
    assert SOL = '1' report "Error in test case #1182/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1183/2803" severity error;
    assert SOR = '0' report "Error in test case #1183/2803" severity error;
    assert SOL = '0' report "Error in test case #1183/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1184/2803" severity error;
    assert SOR = '1' report "Error in test case #1184/2803" severity error;
    assert SOL = '0' report "Error in test case #1184/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1185/2803" severity error;
    assert SOR = '1' report "Error in test case #1185/2803" severity error;
    assert SOL = '0' report "Error in test case #1185/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1186/2803" severity error;
    assert SOR = '1' report "Error in test case #1186/2803" severity error;
    assert SOL = '0' report "Error in test case #1186/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1187/2803" severity error;
    assert SOR = '1' report "Error in test case #1187/2803" severity error;
    assert SOL = '0' report "Error in test case #1187/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1188/2803" severity error;
    assert SOR = '1' report "Error in test case #1188/2803" severity error;
    assert SOL = '0' report "Error in test case #1188/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1189/2803" severity error;
    assert SOR = '1' report "Error in test case #1189/2803" severity error;
    assert SOL = '0' report "Error in test case #1189/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1190/2803" severity error;
    assert SOR = '1' report "Error in test case #1190/2803" severity error;
    assert SOL = '0' report "Error in test case #1190/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1191/2803" severity error;
    assert SOR = '1' report "Error in test case #1191/2803" severity error;
    assert SOL = '0' report "Error in test case #1191/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1192/2803" severity error;
    assert SOR = '0' report "Error in test case #1192/2803" severity error;
    assert SOL = '0' report "Error in test case #1192/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1193/2803" severity error;
    assert SOR = '0' report "Error in test case #1193/2803" severity error;
    assert SOL = '0' report "Error in test case #1193/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1194/2803" severity error;
    assert SOR = '0' report "Error in test case #1194/2803" severity error;
    assert SOL = '0' report "Error in test case #1194/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1195/2803" severity error;
    assert SOR = '0' report "Error in test case #1195/2803" severity error;
    assert SOL = '0' report "Error in test case #1195/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1196/2803" severity error;
    assert SOR = '0' report "Error in test case #1196/2803" severity error;
    assert SOL = '0' report "Error in test case #1196/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1197/2803" severity error;
    assert SOR = '0' report "Error in test case #1197/2803" severity error;
    assert SOL = '0' report "Error in test case #1197/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1198/2803" severity error;
    assert SOR = '0' report "Error in test case #1198/2803" severity error;
    assert SOL = '0' report "Error in test case #1198/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1199/2803" severity error;
    assert SOR = '0' report "Error in test case #1199/2803" severity error;
    assert SOL = '0' report "Error in test case #1199/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1200/2803" severity error;
    assert SOR = '0' report "Error in test case #1200/2803" severity error;
    assert SOL = '0' report "Error in test case #1200/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1201/2803" severity error;
    assert SOR = '0' report "Error in test case #1201/2803" severity error;
    assert SOL = '0' report "Error in test case #1201/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1202/2803" severity error;
    assert SOR = '0' report "Error in test case #1202/2803" severity error;
    assert SOL = '0' report "Error in test case #1202/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "010";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1203/2803" severity error;
    assert SOR = '0' report "Error in test case #1203/2803" severity error;
    assert SOL = '0' report "Error in test case #1203/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1204/2803" severity error;
    assert SOR = '0' report "Error in test case #1204/2803" severity error;
    assert SOL = '0' report "Error in test case #1204/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1205/2803" severity error;
    assert SOR = '0' report "Error in test case #1205/2803" severity error;
    assert SOL = '0' report "Error in test case #1205/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1206/2803" severity error;
    assert SOR = '0' report "Error in test case #1206/2803" severity error;
    assert SOL = '0' report "Error in test case #1206/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1207/2803" severity error;
    assert SOR = '0' report "Error in test case #1207/2803" severity error;
    assert SOL = '0' report "Error in test case #1207/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1208/2803" severity error;
    assert SOR = '0' report "Error in test case #1208/2803" severity error;
    assert SOL = '0' report "Error in test case #1208/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1209/2803" severity error;
    assert SOR = '0' report "Error in test case #1209/2803" severity error;
    assert SOL = '0' report "Error in test case #1209/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1210/2803" severity error;
    assert SOR = '0' report "Error in test case #1210/2803" severity error;
    assert SOL = '0' report "Error in test case #1210/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1211/2803" severity error;
    assert SOR = '0' report "Error in test case #1211/2803" severity error;
    assert SOL = '0' report "Error in test case #1211/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1212/2803" severity error;
    assert SOR = '0' report "Error in test case #1212/2803" severity error;
    assert SOL = '0' report "Error in test case #1212/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1213/2803" severity error;
    assert SOR = '0' report "Error in test case #1213/2803" severity error;
    assert SOL = '0' report "Error in test case #1213/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1214/2803" severity error;
    assert SOR = '0' report "Error in test case #1214/2803" severity error;
    assert SOL = '0' report "Error in test case #1214/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1215/2803" severity error;
    assert SOR = '0' report "Error in test case #1215/2803" severity error;
    assert SOL = '0' report "Error in test case #1215/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1216/2803" severity error;
    assert SOR = '0' report "Error in test case #1216/2803" severity error;
    assert SOL = '0' report "Error in test case #1216/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1217/2803" severity error;
    assert SOR = '0' report "Error in test case #1217/2803" severity error;
    assert SOL = '0' report "Error in test case #1217/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1218/2803" severity error;
    assert SOR = '0' report "Error in test case #1218/2803" severity error;
    assert SOL = '0' report "Error in test case #1218/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1219/2803" severity error;
    assert SOR = '1' report "Error in test case #1219/2803" severity error;
    assert SOL = '1' report "Error in test case #1219/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1220/2803" severity error;
    assert SOR = '1' report "Error in test case #1220/2803" severity error;
    assert SOL = '1' report "Error in test case #1220/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1221/2803" severity error;
    assert SOR = '1' report "Error in test case #1221/2803" severity error;
    assert SOL = '1' report "Error in test case #1221/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1222/2803" severity error;
    assert SOR = '1' report "Error in test case #1222/2803" severity error;
    assert SOL = '1' report "Error in test case #1222/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1223/2803" severity error;
    assert SOR = '1' report "Error in test case #1223/2803" severity error;
    assert SOL = '1' report "Error in test case #1223/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1224/2803" severity error;
    assert SOR = '1' report "Error in test case #1224/2803" severity error;
    assert SOL = '0' report "Error in test case #1224/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1225/2803" severity error;
    assert SOR = '1' report "Error in test case #1225/2803" severity error;
    assert SOL = '0' report "Error in test case #1225/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1226/2803" severity error;
    assert SOR = '1' report "Error in test case #1226/2803" severity error;
    assert SOL = '0' report "Error in test case #1226/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1227/2803" severity error;
    assert SOR = '1' report "Error in test case #1227/2803" severity error;
    assert SOL = '0' report "Error in test case #1227/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1228/2803" severity error;
    assert SOR = '1' report "Error in test case #1228/2803" severity error;
    assert SOL = '0' report "Error in test case #1228/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1229/2803" severity error;
    assert SOR = '1' report "Error in test case #1229/2803" severity error;
    assert SOL = '0' report "Error in test case #1229/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1230/2803" severity error;
    assert SOR = '1' report "Error in test case #1230/2803" severity error;
    assert SOL = '0' report "Error in test case #1230/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1231/2803" severity error;
    assert SOR = '1' report "Error in test case #1231/2803" severity error;
    assert SOL = '0' report "Error in test case #1231/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1232/2803" severity error;
    assert SOR = '0' report "Error in test case #1232/2803" severity error;
    assert SOL = '0' report "Error in test case #1232/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1233/2803" severity error;
    assert SOR = '0' report "Error in test case #1233/2803" severity error;
    assert SOL = '0' report "Error in test case #1233/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1234/2803" severity error;
    assert SOR = '0' report "Error in test case #1234/2803" severity error;
    assert SOL = '0' report "Error in test case #1234/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1235/2803" severity error;
    assert SOR = '0' report "Error in test case #1235/2803" severity error;
    assert SOL = '0' report "Error in test case #1235/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1236/2803" severity error;
    assert SOR = '0' report "Error in test case #1236/2803" severity error;
    assert SOL = '0' report "Error in test case #1236/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1237/2803" severity error;
    assert SOR = '0' report "Error in test case #1237/2803" severity error;
    assert SOL = '0' report "Error in test case #1237/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1238/2803" severity error;
    assert SOR = '0' report "Error in test case #1238/2803" severity error;
    assert SOL = '0' report "Error in test case #1238/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1239/2803" severity error;
    assert SOR = '0' report "Error in test case #1239/2803" severity error;
    assert SOL = '0' report "Error in test case #1239/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1240/2803" severity error;
    assert SOR = '0' report "Error in test case #1240/2803" severity error;
    assert SOL = '0' report "Error in test case #1240/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1241/2803" severity error;
    assert SOR = '0' report "Error in test case #1241/2803" severity error;
    assert SOL = '0' report "Error in test case #1241/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1242/2803" severity error;
    assert SOR = '0' report "Error in test case #1242/2803" severity error;
    assert SOL = '0' report "Error in test case #1242/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1243/2803" severity error;
    assert SOR = '0' report "Error in test case #1243/2803" severity error;
    assert SOL = '0' report "Error in test case #1243/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1244/2803" severity error;
    assert SOR = '0' report "Error in test case #1244/2803" severity error;
    assert SOL = '0' report "Error in test case #1244/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1245/2803" severity error;
    assert SOR = '0' report "Error in test case #1245/2803" severity error;
    assert SOL = '0' report "Error in test case #1245/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1246/2803" severity error;
    assert SOR = '0' report "Error in test case #1246/2803" severity error;
    assert SOL = '0' report "Error in test case #1246/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1247/2803" severity error;
    assert SOR = '0' report "Error in test case #1247/2803" severity error;
    assert SOL = '0' report "Error in test case #1247/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1248/2803" severity error;
    assert SOR = '1' report "Error in test case #1248/2803" severity error;
    assert SOL = '0' report "Error in test case #1248/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1249/2803" severity error;
    assert SOR = '1' report "Error in test case #1249/2803" severity error;
    assert SOL = '0' report "Error in test case #1249/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1250/2803" severity error;
    assert SOR = '1' report "Error in test case #1250/2803" severity error;
    assert SOL = '0' report "Error in test case #1250/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1251/2803" severity error;
    assert SOR = '1' report "Error in test case #1251/2803" severity error;
    assert SOL = '0' report "Error in test case #1251/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1252/2803" severity error;
    assert SOR = '1' report "Error in test case #1252/2803" severity error;
    assert SOL = '0' report "Error in test case #1252/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1253/2803" severity error;
    assert SOR = '1' report "Error in test case #1253/2803" severity error;
    assert SOL = '0' report "Error in test case #1253/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1254/2803" severity error;
    assert SOR = '1' report "Error in test case #1254/2803" severity error;
    assert SOL = '0' report "Error in test case #1254/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1255/2803" severity error;
    assert SOR = '1' report "Error in test case #1255/2803" severity error;
    assert SOL = '0' report "Error in test case #1255/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1256/2803" severity error;
    assert SOR = '1' report "Error in test case #1256/2803" severity error;
    assert SOL = '0' report "Error in test case #1256/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1257/2803" severity error;
    assert SOR = '1' report "Error in test case #1257/2803" severity error;
    assert SOL = '0' report "Error in test case #1257/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1258/2803" severity error;
    assert SOR = '1' report "Error in test case #1258/2803" severity error;
    assert SOL = '0' report "Error in test case #1258/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1259/2803" severity error;
    assert SOR = '1' report "Error in test case #1259/2803" severity error;
    assert SOL = '0' report "Error in test case #1259/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1260/2803" severity error;
    assert SOR = '1' report "Error in test case #1260/2803" severity error;
    assert SOL = '0' report "Error in test case #1260/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1261/2803" severity error;
    assert SOR = '1' report "Error in test case #1261/2803" severity error;
    assert SOL = '0' report "Error in test case #1261/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1262/2803" severity error;
    assert SOR = '1' report "Error in test case #1262/2803" severity error;
    assert SOL = '0' report "Error in test case #1262/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1263/2803" severity error;
    assert SOR = '1' report "Error in test case #1263/2803" severity error;
    assert SOL = '0' report "Error in test case #1263/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1264/2803" severity error;
    assert SOR = '1' report "Error in test case #1264/2803" severity error;
    assert SOL = '0' report "Error in test case #1264/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1265/2803" severity error;
    assert SOR = '1' report "Error in test case #1265/2803" severity error;
    assert SOL = '0' report "Error in test case #1265/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1266/2803" severity error;
    assert SOR = '1' report "Error in test case #1266/2803" severity error;
    assert SOL = '0' report "Error in test case #1266/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1267/2803" severity error;
    assert SOR = '1' report "Error in test case #1267/2803" severity error;
    assert SOL = '0' report "Error in test case #1267/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1268/2803" severity error;
    assert SOR = '1' report "Error in test case #1268/2803" severity error;
    assert SOL = '0' report "Error in test case #1268/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1269/2803" severity error;
    assert SOR = '1' report "Error in test case #1269/2803" severity error;
    assert SOL = '0' report "Error in test case #1269/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1270/2803" severity error;
    assert SOR = '1' report "Error in test case #1270/2803" severity error;
    assert SOL = '0' report "Error in test case #1270/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1271/2803" severity error;
    assert SOR = '1' report "Error in test case #1271/2803" severity error;
    assert SOL = '0' report "Error in test case #1271/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1272/2803" severity error;
    assert SOR = '1' report "Error in test case #1272/2803" severity error;
    assert SOL = '0' report "Error in test case #1272/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1273/2803" severity error;
    assert SOR = '1' report "Error in test case #1273/2803" severity error;
    assert SOL = '0' report "Error in test case #1273/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1274/2803" severity error;
    assert SOR = '1' report "Error in test case #1274/2803" severity error;
    assert SOL = '0' report "Error in test case #1274/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1275/2803" severity error;
    assert SOR = '1' report "Error in test case #1275/2803" severity error;
    assert SOL = '0' report "Error in test case #1275/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1276/2803" severity error;
    assert SOR = '1' report "Error in test case #1276/2803" severity error;
    assert SOL = '0' report "Error in test case #1276/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1277/2803" severity error;
    assert SOR = '1' report "Error in test case #1277/2803" severity error;
    assert SOL = '0' report "Error in test case #1277/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1278/2803" severity error;
    assert SOR = '1' report "Error in test case #1278/2803" severity error;
    assert SOL = '0' report "Error in test case #1278/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000111" report "Error in test case #1279/2803" severity error;
    assert SOR = '1' report "Error in test case #1279/2803" severity error;
    assert SOL = '0' report "Error in test case #1279/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1280/2803" severity error;
    assert SOR = '0' report "Error in test case #1280/2803" severity error;
    assert SOL = '0' report "Error in test case #1280/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1281/2803" severity error;
    assert SOR = '0' report "Error in test case #1281/2803" severity error;
    assert SOL = '0' report "Error in test case #1281/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1282/2803" severity error;
    assert SOR = '0' report "Error in test case #1282/2803" severity error;
    assert SOL = '0' report "Error in test case #1282/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1283/2803" severity error;
    assert SOR = '0' report "Error in test case #1283/2803" severity error;
    assert SOL = '0' report "Error in test case #1283/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1284/2803" severity error;
    assert SOR = '0' report "Error in test case #1284/2803" severity error;
    assert SOL = '0' report "Error in test case #1284/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1285/2803" severity error;
    assert SOR = '0' report "Error in test case #1285/2803" severity error;
    assert SOL = '0' report "Error in test case #1285/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1286/2803" severity error;
    assert SOR = '0' report "Error in test case #1286/2803" severity error;
    assert SOL = '0' report "Error in test case #1286/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1287/2803" severity error;
    assert SOR = '0' report "Error in test case #1287/2803" severity error;
    assert SOL = '0' report "Error in test case #1287/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1288/2803" severity error;
    assert SOR = '0' report "Error in test case #1288/2803" severity error;
    assert SOL = '0' report "Error in test case #1288/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1289/2803" severity error;
    assert SOR = '0' report "Error in test case #1289/2803" severity error;
    assert SOL = '0' report "Error in test case #1289/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1290/2803" severity error;
    assert SOR = '0' report "Error in test case #1290/2803" severity error;
    assert SOL = '0' report "Error in test case #1290/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1291/2803" severity error;
    assert SOR = '0' report "Error in test case #1291/2803" severity error;
    assert SOL = '0' report "Error in test case #1291/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1292/2803" severity error;
    assert SOR = '0' report "Error in test case #1292/2803" severity error;
    assert SOL = '0' report "Error in test case #1292/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1293/2803" severity error;
    assert SOR = '0' report "Error in test case #1293/2803" severity error;
    assert SOL = '0' report "Error in test case #1293/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1294/2803" severity error;
    assert SOR = '0' report "Error in test case #1294/2803" severity error;
    assert SOL = '0' report "Error in test case #1294/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1295/2803" severity error;
    assert SOR = '0' report "Error in test case #1295/2803" severity error;
    assert SOL = '0' report "Error in test case #1295/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1296/2803" severity error;
    assert SOR = '0' report "Error in test case #1296/2803" severity error;
    assert SOL = '0' report "Error in test case #1296/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1297/2803" severity error;
    assert SOR = '0' report "Error in test case #1297/2803" severity error;
    assert SOL = '0' report "Error in test case #1297/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1298/2803" severity error;
    assert SOR = '0' report "Error in test case #1298/2803" severity error;
    assert SOL = '0' report "Error in test case #1298/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1299/2803" severity error;
    assert SOR = '0' report "Error in test case #1299/2803" severity error;
    assert SOL = '0' report "Error in test case #1299/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1300/2803" severity error;
    assert SOR = '0' report "Error in test case #1300/2803" severity error;
    assert SOL = '0' report "Error in test case #1300/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1301/2803" severity error;
    assert SOR = '0' report "Error in test case #1301/2803" severity error;
    assert SOL = '0' report "Error in test case #1301/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1302/2803" severity error;
    assert SOR = '0' report "Error in test case #1302/2803" severity error;
    assert SOL = '0' report "Error in test case #1302/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1303/2803" severity error;
    assert SOR = '0' report "Error in test case #1303/2803" severity error;
    assert SOL = '0' report "Error in test case #1303/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1304/2803" severity error;
    assert SOR = '1' report "Error in test case #1304/2803" severity error;
    assert SOL = '0' report "Error in test case #1304/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1305/2803" severity error;
    assert SOR = '1' report "Error in test case #1305/2803" severity error;
    assert SOL = '0' report "Error in test case #1305/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1306/2803" severity error;
    assert SOR = '1' report "Error in test case #1306/2803" severity error;
    assert SOL = '0' report "Error in test case #1306/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1307/2803" severity error;
    assert SOR = '1' report "Error in test case #1307/2803" severity error;
    assert SOL = '0' report "Error in test case #1307/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1308/2803" severity error;
    assert SOR = '1' report "Error in test case #1308/2803" severity error;
    assert SOL = '0' report "Error in test case #1308/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1309/2803" severity error;
    assert SOR = '1' report "Error in test case #1309/2803" severity error;
    assert SOL = '0' report "Error in test case #1309/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1310/2803" severity error;
    assert SOR = '1' report "Error in test case #1310/2803" severity error;
    assert SOL = '0' report "Error in test case #1310/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1311/2803" severity error;
    assert SOR = '1' report "Error in test case #1311/2803" severity error;
    assert SOL = '0' report "Error in test case #1311/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1312/2803" severity error;
    assert SOR = '0' report "Error in test case #1312/2803" severity error;
    assert SOL = '0' report "Error in test case #1312/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1313/2803" severity error;
    assert SOR = '0' report "Error in test case #1313/2803" severity error;
    assert SOL = '0' report "Error in test case #1313/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1314/2803" severity error;
    assert SOR = '0' report "Error in test case #1314/2803" severity error;
    assert SOL = '0' report "Error in test case #1314/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1315/2803" severity error;
    assert SOR = '0' report "Error in test case #1315/2803" severity error;
    assert SOL = '0' report "Error in test case #1315/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1316/2803" severity error;
    assert SOR = '0' report "Error in test case #1316/2803" severity error;
    assert SOL = '0' report "Error in test case #1316/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1317/2803" severity error;
    assert SOR = '0' report "Error in test case #1317/2803" severity error;
    assert SOL = '0' report "Error in test case #1317/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1318/2803" severity error;
    assert SOR = '0' report "Error in test case #1318/2803" severity error;
    assert SOL = '0' report "Error in test case #1318/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1319/2803" severity error;
    assert SOR = '0' report "Error in test case #1319/2803" severity error;
    assert SOL = '0' report "Error in test case #1319/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1320/2803" severity error;
    assert SOR = '1' report "Error in test case #1320/2803" severity error;
    assert SOL = '0' report "Error in test case #1320/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1321/2803" severity error;
    assert SOR = '1' report "Error in test case #1321/2803" severity error;
    assert SOL = '0' report "Error in test case #1321/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1322/2803" severity error;
    assert SOR = '1' report "Error in test case #1322/2803" severity error;
    assert SOL = '0' report "Error in test case #1322/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1323/2803" severity error;
    assert SOR = '1' report "Error in test case #1323/2803" severity error;
    assert SOL = '0' report "Error in test case #1323/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1324/2803" severity error;
    assert SOR = '1' report "Error in test case #1324/2803" severity error;
    assert SOL = '0' report "Error in test case #1324/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1325/2803" severity error;
    assert SOR = '0' report "Error in test case #1325/2803" severity error;
    assert SOL = '0' report "Error in test case #1325/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1326/2803" severity error;
    assert SOR = '0' report "Error in test case #1326/2803" severity error;
    assert SOL = '0' report "Error in test case #1326/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1327/2803" severity error;
    assert SOR = '0' report "Error in test case #1327/2803" severity error;
    assert SOL = '0' report "Error in test case #1327/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1328/2803" severity error;
    assert SOR = '1' report "Error in test case #1328/2803" severity error;
    assert SOL = '0' report "Error in test case #1328/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1329/2803" severity error;
    assert SOR = '1' report "Error in test case #1329/2803" severity error;
    assert SOL = '0' report "Error in test case #1329/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1330/2803" severity error;
    assert SOR = '1' report "Error in test case #1330/2803" severity error;
    assert SOL = '0' report "Error in test case #1330/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1331/2803" severity error;
    assert SOR = '1' report "Error in test case #1331/2803" severity error;
    assert SOL = '0' report "Error in test case #1331/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1332/2803" severity error;
    assert SOR = '1' report "Error in test case #1332/2803" severity error;
    assert SOL = '0' report "Error in test case #1332/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1333/2803" severity error;
    assert SOR = '1' report "Error in test case #1333/2803" severity error;
    assert SOL = '0' report "Error in test case #1333/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1334/2803" severity error;
    assert SOR = '1' report "Error in test case #1334/2803" severity error;
    assert SOL = '0' report "Error in test case #1334/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1335/2803" severity error;
    assert SOR = '1' report "Error in test case #1335/2803" severity error;
    assert SOL = '0' report "Error in test case #1335/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1336/2803" severity error;
    assert SOR = '0' report "Error in test case #1336/2803" severity error;
    assert SOL = '0' report "Error in test case #1336/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1337/2803" severity error;
    assert SOR = '0' report "Error in test case #1337/2803" severity error;
    assert SOL = '0' report "Error in test case #1337/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1338/2803" severity error;
    assert SOR = '0' report "Error in test case #1338/2803" severity error;
    assert SOL = '0' report "Error in test case #1338/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1339/2803" severity error;
    assert SOR = '0' report "Error in test case #1339/2803" severity error;
    assert SOL = '0' report "Error in test case #1339/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1340/2803" severity error;
    assert SOR = '0' report "Error in test case #1340/2803" severity error;
    assert SOL = '0' report "Error in test case #1340/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1341/2803" severity error;
    assert SOR = '0' report "Error in test case #1341/2803" severity error;
    assert SOL = '0' report "Error in test case #1341/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1342/2803" severity error;
    assert SOR = '0' report "Error in test case #1342/2803" severity error;
    assert SOL = '0' report "Error in test case #1342/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1343/2803" severity error;
    assert SOR = '0' report "Error in test case #1343/2803" severity error;
    assert SOL = '0' report "Error in test case #1343/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1344/2803" severity error;
    assert SOR = '0' report "Error in test case #1344/2803" severity error;
    assert SOL = '0' report "Error in test case #1344/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1345/2803" severity error;
    assert SOR = '0' report "Error in test case #1345/2803" severity error;
    assert SOL = '0' report "Error in test case #1345/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1346/2803" severity error;
    assert SOR = '0' report "Error in test case #1346/2803" severity error;
    assert SOL = '0' report "Error in test case #1346/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1347/2803" severity error;
    assert SOR = '0' report "Error in test case #1347/2803" severity error;
    assert SOL = '0' report "Error in test case #1347/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1348/2803" severity error;
    assert SOR = '0' report "Error in test case #1348/2803" severity error;
    assert SOL = '0' report "Error in test case #1348/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1349/2803" severity error;
    assert SOR = '0' report "Error in test case #1349/2803" severity error;
    assert SOL = '0' report "Error in test case #1349/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1350/2803" severity error;
    assert SOR = '0' report "Error in test case #1350/2803" severity error;
    assert SOL = '0' report "Error in test case #1350/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1351/2803" severity error;
    assert SOR = '0' report "Error in test case #1351/2803" severity error;
    assert SOL = '0' report "Error in test case #1351/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1352/2803" severity error;
    assert SOR = '0' report "Error in test case #1352/2803" severity error;
    assert SOL = '0' report "Error in test case #1352/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1353/2803" severity error;
    assert SOR = '0' report "Error in test case #1353/2803" severity error;
    assert SOL = '0' report "Error in test case #1353/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1354/2803" severity error;
    assert SOR = '0' report "Error in test case #1354/2803" severity error;
    assert SOL = '0' report "Error in test case #1354/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1355/2803" severity error;
    assert SOR = '0' report "Error in test case #1355/2803" severity error;
    assert SOL = '0' report "Error in test case #1355/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1356/2803" severity error;
    assert SOR = '0' report "Error in test case #1356/2803" severity error;
    assert SOL = '0' report "Error in test case #1356/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1357/2803" severity error;
    assert SOR = '0' report "Error in test case #1357/2803" severity error;
    assert SOL = '0' report "Error in test case #1357/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1358/2803" severity error;
    assert SOR = '0' report "Error in test case #1358/2803" severity error;
    assert SOL = '0' report "Error in test case #1358/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1359/2803" severity error;
    assert SOR = '0' report "Error in test case #1359/2803" severity error;
    assert SOL = '0' report "Error in test case #1359/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1360/2803" severity error;
    assert SOR = '1' report "Error in test case #1360/2803" severity error;
    assert SOL = '0' report "Error in test case #1360/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1361/2803" severity error;
    assert SOR = '1' report "Error in test case #1361/2803" severity error;
    assert SOL = '0' report "Error in test case #1361/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1362/2803" severity error;
    assert SOR = '1' report "Error in test case #1362/2803" severity error;
    assert SOL = '0' report "Error in test case #1362/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1363/2803" severity error;
    assert SOR = '1' report "Error in test case #1363/2803" severity error;
    assert SOL = '0' report "Error in test case #1363/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1364/2803" severity error;
    assert SOR = '1' report "Error in test case #1364/2803" severity error;
    assert SOL = '0' report "Error in test case #1364/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1365/2803" severity error;
    assert SOR = '1' report "Error in test case #1365/2803" severity error;
    assert SOL = '0' report "Error in test case #1365/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1366/2803" severity error;
    assert SOR = '1' report "Error in test case #1366/2803" severity error;
    assert SOL = '0' report "Error in test case #1366/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1367/2803" severity error;
    assert SOR = '1' report "Error in test case #1367/2803" severity error;
    assert SOL = '0' report "Error in test case #1367/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1368/2803" severity error;
    assert SOR = '0' report "Error in test case #1368/2803" severity error;
    assert SOL = '0' report "Error in test case #1368/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1369/2803" severity error;
    assert SOR = '0' report "Error in test case #1369/2803" severity error;
    assert SOL = '0' report "Error in test case #1369/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1370/2803" severity error;
    assert SOR = '0' report "Error in test case #1370/2803" severity error;
    assert SOL = '0' report "Error in test case #1370/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1371/2803" severity error;
    assert SOR = '0' report "Error in test case #1371/2803" severity error;
    assert SOL = '0' report "Error in test case #1371/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1372/2803" severity error;
    assert SOR = '0' report "Error in test case #1372/2803" severity error;
    assert SOL = '0' report "Error in test case #1372/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1373/2803" severity error;
    assert SOR = '0' report "Error in test case #1373/2803" severity error;
    assert SOL = '0' report "Error in test case #1373/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1374/2803" severity error;
    assert SOR = '0' report "Error in test case #1374/2803" severity error;
    assert SOL = '0' report "Error in test case #1374/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1375/2803" severity error;
    assert SOR = '0' report "Error in test case #1375/2803" severity error;
    assert SOL = '0' report "Error in test case #1375/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1376/2803" severity error;
    assert SOR = '0' report "Error in test case #1376/2803" severity error;
    assert SOL = '0' report "Error in test case #1376/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1377/2803" severity error;
    assert SOR = '0' report "Error in test case #1377/2803" severity error;
    assert SOL = '0' report "Error in test case #1377/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1378/2803" severity error;
    assert SOR = '0' report "Error in test case #1378/2803" severity error;
    assert SOL = '0' report "Error in test case #1378/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1379/2803" severity error;
    assert SOR = '0' report "Error in test case #1379/2803" severity error;
    assert SOL = '0' report "Error in test case #1379/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1380/2803" severity error;
    assert SOR = '0' report "Error in test case #1380/2803" severity error;
    assert SOL = '0' report "Error in test case #1380/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1381/2803" severity error;
    assert SOR = '0' report "Error in test case #1381/2803" severity error;
    assert SOL = '0' report "Error in test case #1381/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1382/2803" severity error;
    assert SOR = '0' report "Error in test case #1382/2803" severity error;
    assert SOL = '0' report "Error in test case #1382/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1383/2803" severity error;
    assert SOR = '0' report "Error in test case #1383/2803" severity error;
    assert SOL = '0' report "Error in test case #1383/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1384/2803" severity error;
    assert SOR = '0' report "Error in test case #1384/2803" severity error;
    assert SOL = '0' report "Error in test case #1384/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1385/2803" severity error;
    assert SOR = '0' report "Error in test case #1385/2803" severity error;
    assert SOL = '0' report "Error in test case #1385/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1386/2803" severity error;
    assert SOR = '0' report "Error in test case #1386/2803" severity error;
    assert SOL = '0' report "Error in test case #1386/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1387/2803" severity error;
    assert SOR = '0' report "Error in test case #1387/2803" severity error;
    assert SOL = '0' report "Error in test case #1387/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1388/2803" severity error;
    assert SOR = '0' report "Error in test case #1388/2803" severity error;
    assert SOL = '0' report "Error in test case #1388/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1389/2803" severity error;
    assert SOR = '0' report "Error in test case #1389/2803" severity error;
    assert SOL = '0' report "Error in test case #1389/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1390/2803" severity error;
    assert SOR = '0' report "Error in test case #1390/2803" severity error;
    assert SOL = '0' report "Error in test case #1390/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1391/2803" severity error;
    assert SOR = '0' report "Error in test case #1391/2803" severity error;
    assert SOL = '0' report "Error in test case #1391/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1392/2803" severity error;
    assert SOR = '0' report "Error in test case #1392/2803" severity error;
    assert SOL = '0' report "Error in test case #1392/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1393/2803" severity error;
    assert SOR = '0' report "Error in test case #1393/2803" severity error;
    assert SOL = '0' report "Error in test case #1393/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1394/2803" severity error;
    assert SOR = '0' report "Error in test case #1394/2803" severity error;
    assert SOL = '0' report "Error in test case #1394/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1395/2803" severity error;
    assert SOR = '0' report "Error in test case #1395/2803" severity error;
    assert SOL = '0' report "Error in test case #1395/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1396/2803" severity error;
    assert SOR = '0' report "Error in test case #1396/2803" severity error;
    assert SOL = '0' report "Error in test case #1396/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1397/2803" severity error;
    assert SOR = '0' report "Error in test case #1397/2803" severity error;
    assert SOL = '0' report "Error in test case #1397/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1398/2803" severity error;
    assert SOR = '0' report "Error in test case #1398/2803" severity error;
    assert SOL = '0' report "Error in test case #1398/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1399/2803" severity error;
    assert SOR = '0' report "Error in test case #1399/2803" severity error;
    assert SOL = '0' report "Error in test case #1399/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1400/2803" severity error;
    assert SOR = '1' report "Error in test case #1400/2803" severity error;
    assert SOL = '0' report "Error in test case #1400/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1401/2803" severity error;
    assert SOR = '1' report "Error in test case #1401/2803" severity error;
    assert SOL = '0' report "Error in test case #1401/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1402/2803" severity error;
    assert SOR = '1' report "Error in test case #1402/2803" severity error;
    assert SOL = '0' report "Error in test case #1402/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1403/2803" severity error;
    assert SOR = '1' report "Error in test case #1403/2803" severity error;
    assert SOL = '0' report "Error in test case #1403/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1404/2803" severity error;
    assert SOR = '1' report "Error in test case #1404/2803" severity error;
    assert SOL = '0' report "Error in test case #1404/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1405/2803" severity error;
    assert SOR = '1' report "Error in test case #1405/2803" severity error;
    assert SOL = '0' report "Error in test case #1405/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1406/2803" severity error;
    assert SOR = '1' report "Error in test case #1406/2803" severity error;
    assert SOL = '0' report "Error in test case #1406/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1407/2803" severity error;
    assert SOR = '1' report "Error in test case #1407/2803" severity error;
    assert SOL = '0' report "Error in test case #1407/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1408/2803" severity error;
    assert SOR = '0' report "Error in test case #1408/2803" severity error;
    assert SOL = '0' report "Error in test case #1408/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1409/2803" severity error;
    assert SOR = '0' report "Error in test case #1409/2803" severity error;
    assert SOL = '0' report "Error in test case #1409/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1410/2803" severity error;
    assert SOR = '0' report "Error in test case #1410/2803" severity error;
    assert SOL = '0' report "Error in test case #1410/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1411/2803" severity error;
    assert SOR = '0' report "Error in test case #1411/2803" severity error;
    assert SOL = '0' report "Error in test case #1411/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1412/2803" severity error;
    assert SOR = '0' report "Error in test case #1412/2803" severity error;
    assert SOL = '0' report "Error in test case #1412/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1413/2803" severity error;
    assert SOR = '0' report "Error in test case #1413/2803" severity error;
    assert SOL = '0' report "Error in test case #1413/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1414/2803" severity error;
    assert SOR = '0' report "Error in test case #1414/2803" severity error;
    assert SOL = '0' report "Error in test case #1414/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1415/2803" severity error;
    assert SOR = '0' report "Error in test case #1415/2803" severity error;
    assert SOL = '0' report "Error in test case #1415/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1416/2803" severity error;
    assert SOR = '0' report "Error in test case #1416/2803" severity error;
    assert SOL = '0' report "Error in test case #1416/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1417/2803" severity error;
    assert SOR = '0' report "Error in test case #1417/2803" severity error;
    assert SOL = '0' report "Error in test case #1417/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1418/2803" severity error;
    assert SOR = '0' report "Error in test case #1418/2803" severity error;
    assert SOL = '0' report "Error in test case #1418/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1419/2803" severity error;
    assert SOR = '0' report "Error in test case #1419/2803" severity error;
    assert SOL = '0' report "Error in test case #1419/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1420/2803" severity error;
    assert SOR = '0' report "Error in test case #1420/2803" severity error;
    assert SOL = '0' report "Error in test case #1420/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1421/2803" severity error;
    assert SOR = '0' report "Error in test case #1421/2803" severity error;
    assert SOL = '0' report "Error in test case #1421/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1422/2803" severity error;
    assert SOR = '0' report "Error in test case #1422/2803" severity error;
    assert SOL = '0' report "Error in test case #1422/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1423/2803" severity error;
    assert SOR = '0' report "Error in test case #1423/2803" severity error;
    assert SOL = '0' report "Error in test case #1423/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1424/2803" severity error;
    assert SOR = '0' report "Error in test case #1424/2803" severity error;
    assert SOL = '0' report "Error in test case #1424/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1425/2803" severity error;
    assert SOR = '0' report "Error in test case #1425/2803" severity error;
    assert SOL = '0' report "Error in test case #1425/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1426/2803" severity error;
    assert SOR = '0' report "Error in test case #1426/2803" severity error;
    assert SOL = '0' report "Error in test case #1426/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1427/2803" severity error;
    assert SOR = '0' report "Error in test case #1427/2803" severity error;
    assert SOL = '0' report "Error in test case #1427/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1428/2803" severity error;
    assert SOR = '0' report "Error in test case #1428/2803" severity error;
    assert SOL = '0' report "Error in test case #1428/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1429/2803" severity error;
    assert SOR = '0' report "Error in test case #1429/2803" severity error;
    assert SOL = '0' report "Error in test case #1429/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1430/2803" severity error;
    assert SOR = '0' report "Error in test case #1430/2803" severity error;
    assert SOL = '0' report "Error in test case #1430/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1431/2803" severity error;
    assert SOR = '0' report "Error in test case #1431/2803" severity error;
    assert SOL = '0' report "Error in test case #1431/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1432/2803" severity error;
    assert SOR = '0' report "Error in test case #1432/2803" severity error;
    assert SOL = '0' report "Error in test case #1432/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1433/2803" severity error;
    assert SOR = '0' report "Error in test case #1433/2803" severity error;
    assert SOL = '0' report "Error in test case #1433/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1434/2803" severity error;
    assert SOR = '0' report "Error in test case #1434/2803" severity error;
    assert SOL = '0' report "Error in test case #1434/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1435/2803" severity error;
    assert SOR = '0' report "Error in test case #1435/2803" severity error;
    assert SOL = '0' report "Error in test case #1435/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1436/2803" severity error;
    assert SOR = '1' report "Error in test case #1436/2803" severity error;
    assert SOL = '1' report "Error in test case #1436/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1437/2803" severity error;
    assert SOR = '1' report "Error in test case #1437/2803" severity error;
    assert SOL = '1' report "Error in test case #1437/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1438/2803" severity error;
    assert SOR = '1' report "Error in test case #1438/2803" severity error;
    assert SOL = '1' report "Error in test case #1438/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1439/2803" severity error;
    assert SOR = '1' report "Error in test case #1439/2803" severity error;
    assert SOL = '1' report "Error in test case #1439/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1440/2803" severity error;
    assert SOR = '0' report "Error in test case #1440/2803" severity error;
    assert SOL = '0' report "Error in test case #1440/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1441/2803" severity error;
    assert SOR = '0' report "Error in test case #1441/2803" severity error;
    assert SOL = '0' report "Error in test case #1441/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1442/2803" severity error;
    assert SOR = '0' report "Error in test case #1442/2803" severity error;
    assert SOL = '0' report "Error in test case #1442/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1443/2803" severity error;
    assert SOR = '0' report "Error in test case #1443/2803" severity error;
    assert SOL = '0' report "Error in test case #1443/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1444/2803" severity error;
    assert SOR = '0' report "Error in test case #1444/2803" severity error;
    assert SOL = '0' report "Error in test case #1444/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1445/2803" severity error;
    assert SOR = '0' report "Error in test case #1445/2803" severity error;
    assert SOL = '0' report "Error in test case #1445/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1446/2803" severity error;
    assert SOR = '0' report "Error in test case #1446/2803" severity error;
    assert SOL = '0' report "Error in test case #1446/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1447/2803" severity error;
    assert SOR = '0' report "Error in test case #1447/2803" severity error;
    assert SOL = '0' report "Error in test case #1447/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1448/2803" severity error;
    assert SOR = '0' report "Error in test case #1448/2803" severity error;
    assert SOL = '0' report "Error in test case #1448/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1449/2803" severity error;
    assert SOR = '0' report "Error in test case #1449/2803" severity error;
    assert SOL = '0' report "Error in test case #1449/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1450/2803" severity error;
    assert SOR = '0' report "Error in test case #1450/2803" severity error;
    assert SOL = '0' report "Error in test case #1450/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1451/2803" severity error;
    assert SOR = '0' report "Error in test case #1451/2803" severity error;
    assert SOL = '0' report "Error in test case #1451/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1452/2803" severity error;
    assert SOR = '0' report "Error in test case #1452/2803" severity error;
    assert SOL = '0' report "Error in test case #1452/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1453/2803" severity error;
    assert SOR = '0' report "Error in test case #1453/2803" severity error;
    assert SOL = '0' report "Error in test case #1453/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1454/2803" severity error;
    assert SOR = '0' report "Error in test case #1454/2803" severity error;
    assert SOL = '0' report "Error in test case #1454/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1455/2803" severity error;
    assert SOR = '0' report "Error in test case #1455/2803" severity error;
    assert SOL = '0' report "Error in test case #1455/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1456/2803" severity error;
    assert SOR = '1' report "Error in test case #1456/2803" severity error;
    assert SOL = '0' report "Error in test case #1456/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1457/2803" severity error;
    assert SOR = '1' report "Error in test case #1457/2803" severity error;
    assert SOL = '0' report "Error in test case #1457/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1458/2803" severity error;
    assert SOR = '1' report "Error in test case #1458/2803" severity error;
    assert SOL = '0' report "Error in test case #1458/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1459/2803" severity error;
    assert SOR = '1' report "Error in test case #1459/2803" severity error;
    assert SOL = '0' report "Error in test case #1459/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1460/2803" severity error;
    assert SOR = '1' report "Error in test case #1460/2803" severity error;
    assert SOL = '0' report "Error in test case #1460/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1461/2803" severity error;
    assert SOR = '1' report "Error in test case #1461/2803" severity error;
    assert SOL = '0' report "Error in test case #1461/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1462/2803" severity error;
    assert SOR = '1' report "Error in test case #1462/2803" severity error;
    assert SOL = '0' report "Error in test case #1462/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1463/2803" severity error;
    assert SOR = '1' report "Error in test case #1463/2803" severity error;
    assert SOL = '0' report "Error in test case #1463/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1464/2803" severity error;
    assert SOR = '0' report "Error in test case #1464/2803" severity error;
    assert SOL = '0' report "Error in test case #1464/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1465/2803" severity error;
    assert SOR = '0' report "Error in test case #1465/2803" severity error;
    assert SOL = '0' report "Error in test case #1465/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1466/2803" severity error;
    assert SOR = '0' report "Error in test case #1466/2803" severity error;
    assert SOL = '0' report "Error in test case #1466/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1467/2803" severity error;
    assert SOR = '0' report "Error in test case #1467/2803" severity error;
    assert SOL = '0' report "Error in test case #1467/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1468/2803" severity error;
    assert SOR = '0' report "Error in test case #1468/2803" severity error;
    assert SOL = '0' report "Error in test case #1468/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1469/2803" severity error;
    assert SOR = '0' report "Error in test case #1469/2803" severity error;
    assert SOL = '0' report "Error in test case #1469/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1470/2803" severity error;
    assert SOR = '0' report "Error in test case #1470/2803" severity error;
    assert SOL = '0' report "Error in test case #1470/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1471/2803" severity error;
    assert SOR = '0' report "Error in test case #1471/2803" severity error;
    assert SOL = '0' report "Error in test case #1471/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1472/2803" severity error;
    assert SOR = '0' report "Error in test case #1472/2803" severity error;
    assert SOL = '0' report "Error in test case #1472/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1473/2803" severity error;
    assert SOR = '0' report "Error in test case #1473/2803" severity error;
    assert SOL = '0' report "Error in test case #1473/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1474/2803" severity error;
    assert SOR = '0' report "Error in test case #1474/2803" severity error;
    assert SOL = '0' report "Error in test case #1474/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1475/2803" severity error;
    assert SOR = '0' report "Error in test case #1475/2803" severity error;
    assert SOL = '0' report "Error in test case #1475/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1476/2803" severity error;
    assert SOR = '0' report "Error in test case #1476/2803" severity error;
    assert SOL = '0' report "Error in test case #1476/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1477/2803" severity error;
    assert SOR = '0' report "Error in test case #1477/2803" severity error;
    assert SOL = '0' report "Error in test case #1477/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1478/2803" severity error;
    assert SOR = '0' report "Error in test case #1478/2803" severity error;
    assert SOL = '0' report "Error in test case #1478/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1479/2803" severity error;
    assert SOR = '0' report "Error in test case #1479/2803" severity error;
    assert SOL = '0' report "Error in test case #1479/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1480/2803" severity error;
    assert SOR = '0' report "Error in test case #1480/2803" severity error;
    assert SOL = '0' report "Error in test case #1480/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1481/2803" severity error;
    assert SOR = '0' report "Error in test case #1481/2803" severity error;
    assert SOL = '0' report "Error in test case #1481/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1482/2803" severity error;
    assert SOR = '0' report "Error in test case #1482/2803" severity error;
    assert SOL = '0' report "Error in test case #1482/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1483/2803" severity error;
    assert SOR = '0' report "Error in test case #1483/2803" severity error;
    assert SOL = '0' report "Error in test case #1483/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1484/2803" severity error;
    assert SOR = '0' report "Error in test case #1484/2803" severity error;
    assert SOL = '0' report "Error in test case #1484/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1485/2803" severity error;
    assert SOR = '0' report "Error in test case #1485/2803" severity error;
    assert SOL = '0' report "Error in test case #1485/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1486/2803" severity error;
    assert SOR = '0' report "Error in test case #1486/2803" severity error;
    assert SOL = '0' report "Error in test case #1486/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1487/2803" severity error;
    assert SOR = '0' report "Error in test case #1487/2803" severity error;
    assert SOL = '0' report "Error in test case #1487/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1488/2803" severity error;
    assert SOR = '0' report "Error in test case #1488/2803" severity error;
    assert SOL = '0' report "Error in test case #1488/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1489/2803" severity error;
    assert SOR = '0' report "Error in test case #1489/2803" severity error;
    assert SOL = '0' report "Error in test case #1489/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1490/2803" severity error;
    assert SOR = '0' report "Error in test case #1490/2803" severity error;
    assert SOL = '0' report "Error in test case #1490/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1491/2803" severity error;
    assert SOR = '0' report "Error in test case #1491/2803" severity error;
    assert SOL = '0' report "Error in test case #1491/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1492/2803" severity error;
    assert SOR = '1' report "Error in test case #1492/2803" severity error;
    assert SOL = '1' report "Error in test case #1492/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1493/2803" severity error;
    assert SOR = '1' report "Error in test case #1493/2803" severity error;
    assert SOL = '1' report "Error in test case #1493/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1494/2803" severity error;
    assert SOR = '1' report "Error in test case #1494/2803" severity error;
    assert SOL = '1' report "Error in test case #1494/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1495/2803" severity error;
    assert SOR = '1' report "Error in test case #1495/2803" severity error;
    assert SOL = '1' report "Error in test case #1495/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1496/2803" severity error;
    assert SOR = '0' report "Error in test case #1496/2803" severity error;
    assert SOL = '0' report "Error in test case #1496/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1497/2803" severity error;
    assert SOR = '0' report "Error in test case #1497/2803" severity error;
    assert SOL = '0' report "Error in test case #1497/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1498/2803" severity error;
    assert SOR = '0' report "Error in test case #1498/2803" severity error;
    assert SOL = '0' report "Error in test case #1498/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1499/2803" severity error;
    assert SOR = '0' report "Error in test case #1499/2803" severity error;
    assert SOL = '0' report "Error in test case #1499/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1500/2803" severity error;
    assert SOR = '0' report "Error in test case #1500/2803" severity error;
    assert SOL = '0' report "Error in test case #1500/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1501/2803" severity error;
    assert SOR = '0' report "Error in test case #1501/2803" severity error;
    assert SOL = '0' report "Error in test case #1501/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1502/2803" severity error;
    assert SOR = '0' report "Error in test case #1502/2803" severity error;
    assert SOL = '0' report "Error in test case #1502/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1503/2803" severity error;
    assert SOR = '0' report "Error in test case #1503/2803" severity error;
    assert SOL = '0' report "Error in test case #1503/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1504/2803" severity error;
    assert SOR = '0' report "Error in test case #1504/2803" severity error;
    assert SOL = '0' report "Error in test case #1504/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1505/2803" severity error;
    assert SOR = '0' report "Error in test case #1505/2803" severity error;
    assert SOL = '0' report "Error in test case #1505/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1506/2803" severity error;
    assert SOR = '0' report "Error in test case #1506/2803" severity error;
    assert SOL = '0' report "Error in test case #1506/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1507/2803" severity error;
    assert SOR = '0' report "Error in test case #1507/2803" severity error;
    assert SOL = '0' report "Error in test case #1507/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1508/2803" severity error;
    assert SOR = '0' report "Error in test case #1508/2803" severity error;
    assert SOL = '0' report "Error in test case #1508/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1509/2803" severity error;
    assert SOR = '0' report "Error in test case #1509/2803" severity error;
    assert SOL = '0' report "Error in test case #1509/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1510/2803" severity error;
    assert SOR = '0' report "Error in test case #1510/2803" severity error;
    assert SOL = '0' report "Error in test case #1510/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000010" report "Error in test case #1511/2803" severity error;
    assert SOR = '0' report "Error in test case #1511/2803" severity error;
    assert SOL = '0' report "Error in test case #1511/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1512/2803" severity error;
    assert SOR = '1' report "Error in test case #1512/2803" severity error;
    assert SOL = '0' report "Error in test case #1512/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1513/2803" severity error;
    assert SOR = '1' report "Error in test case #1513/2803" severity error;
    assert SOL = '0' report "Error in test case #1513/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1514/2803" severity error;
    assert SOR = '1' report "Error in test case #1514/2803" severity error;
    assert SOL = '0' report "Error in test case #1514/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1515/2803" severity error;
    assert SOR = '1' report "Error in test case #1515/2803" severity error;
    assert SOL = '0' report "Error in test case #1515/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1516/2803" severity error;
    assert SOR = '1' report "Error in test case #1516/2803" severity error;
    assert SOL = '0' report "Error in test case #1516/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1517/2803" severity error;
    assert SOR = '0' report "Error in test case #1517/2803" severity error;
    assert SOL = '0' report "Error in test case #1517/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1518/2803" severity error;
    assert SOR = '0' report "Error in test case #1518/2803" severity error;
    assert SOL = '0' report "Error in test case #1518/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1519/2803" severity error;
    assert SOR = '0' report "Error in test case #1519/2803" severity error;
    assert SOL = '0' report "Error in test case #1519/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1520/2803" severity error;
    assert SOR = '0' report "Error in test case #1520/2803" severity error;
    assert SOL = '0' report "Error in test case #1520/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1521/2803" severity error;
    assert SOR = '0' report "Error in test case #1521/2803" severity error;
    assert SOL = '0' report "Error in test case #1521/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1522/2803" severity error;
    assert SOR = '0' report "Error in test case #1522/2803" severity error;
    assert SOL = '0' report "Error in test case #1522/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1523/2803" severity error;
    assert SOR = '0' report "Error in test case #1523/2803" severity error;
    assert SOL = '0' report "Error in test case #1523/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1524/2803" severity error;
    assert SOR = '0' report "Error in test case #1524/2803" severity error;
    assert SOL = '0' report "Error in test case #1524/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1525/2803" severity error;
    assert SOR = '0' report "Error in test case #1525/2803" severity error;
    assert SOL = '0' report "Error in test case #1525/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1526/2803" severity error;
    assert SOR = '0' report "Error in test case #1526/2803" severity error;
    assert SOL = '0' report "Error in test case #1526/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1527/2803" severity error;
    assert SOR = '0' report "Error in test case #1527/2803" severity error;
    assert SOL = '0' report "Error in test case #1527/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1528/2803" severity error;
    assert SOR = '1' report "Error in test case #1528/2803" severity error;
    assert SOL = '0' report "Error in test case #1528/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1529/2803" severity error;
    assert SOR = '1' report "Error in test case #1529/2803" severity error;
    assert SOL = '0' report "Error in test case #1529/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1530/2803" severity error;
    assert SOR = '1' report "Error in test case #1530/2803" severity error;
    assert SOL = '0' report "Error in test case #1530/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1531/2803" severity error;
    assert SOR = '1' report "Error in test case #1531/2803" severity error;
    assert SOL = '0' report "Error in test case #1531/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1532/2803" severity error;
    assert SOR = '1' report "Error in test case #1532/2803" severity error;
    assert SOL = '0' report "Error in test case #1532/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1533/2803" severity error;
    assert SOR = '0' report "Error in test case #1533/2803" severity error;
    assert SOL = '0' report "Error in test case #1533/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1534/2803" severity error;
    assert SOR = '0' report "Error in test case #1534/2803" severity error;
    assert SOL = '0' report "Error in test case #1534/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1535/2803" severity error;
    assert SOR = '0' report "Error in test case #1535/2803" severity error;
    assert SOL = '0' report "Error in test case #1535/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1536/2803" severity error;
    assert SOR = '0' report "Error in test case #1536/2803" severity error;
    assert SOL = '0' report "Error in test case #1536/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1537/2803" severity error;
    assert SOR = '0' report "Error in test case #1537/2803" severity error;
    assert SOL = '0' report "Error in test case #1537/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1538/2803" severity error;
    assert SOR = '0' report "Error in test case #1538/2803" severity error;
    assert SOL = '0' report "Error in test case #1538/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1539/2803" severity error;
    assert SOR = '0' report "Error in test case #1539/2803" severity error;
    assert SOL = '0' report "Error in test case #1539/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000100" report "Error in test case #1540/2803" severity error;
    assert SOR = '0' report "Error in test case #1540/2803" severity error;
    assert SOL = '0' report "Error in test case #1540/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1541/2803" severity error;
    assert SOR = '0' report "Error in test case #1541/2803" severity error;
    assert SOL = '0' report "Error in test case #1541/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1542/2803" severity error;
    assert SOR = '0' report "Error in test case #1542/2803" severity error;
    assert SOL = '0' report "Error in test case #1542/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1543/2803" severity error;
    assert SOR = '0' report "Error in test case #1543/2803" severity error;
    assert SOL = '0' report "Error in test case #1543/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1544/2803" severity error;
    assert SOR = '1' report "Error in test case #1544/2803" severity error;
    assert SOL = '0' report "Error in test case #1544/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1545/2803" severity error;
    assert SOR = '1' report "Error in test case #1545/2803" severity error;
    assert SOL = '0' report "Error in test case #1545/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1546/2803" severity error;
    assert SOR = '1' report "Error in test case #1546/2803" severity error;
    assert SOL = '0' report "Error in test case #1546/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1547/2803" severity error;
    assert SOR = '1' report "Error in test case #1547/2803" severity error;
    assert SOL = '0' report "Error in test case #1547/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1548/2803" severity error;
    assert SOR = '1' report "Error in test case #1548/2803" severity error;
    assert SOL = '0' report "Error in test case #1548/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1549/2803" severity error;
    assert SOR = '1' report "Error in test case #1549/2803" severity error;
    assert SOL = '0' report "Error in test case #1549/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1550/2803" severity error;
    assert SOR = '1' report "Error in test case #1550/2803" severity error;
    assert SOL = '0' report "Error in test case #1550/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1551/2803" severity error;
    assert SOR = '1' report "Error in test case #1551/2803" severity error;
    assert SOL = '0' report "Error in test case #1551/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1552/2803" severity error;
    assert SOR = '1' report "Error in test case #1552/2803" severity error;
    assert SOL = '0' report "Error in test case #1552/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1553/2803" severity error;
    assert SOR = '1' report "Error in test case #1553/2803" severity error;
    assert SOL = '0' report "Error in test case #1553/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1554/2803" severity error;
    assert SOR = '1' report "Error in test case #1554/2803" severity error;
    assert SOL = '0' report "Error in test case #1554/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1555/2803" severity error;
    assert SOR = '1' report "Error in test case #1555/2803" severity error;
    assert SOL = '0' report "Error in test case #1555/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1556/2803" severity error;
    assert SOR = '1' report "Error in test case #1556/2803" severity error;
    assert SOL = '0' report "Error in test case #1556/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1557/2803" severity error;
    assert SOR = '1' report "Error in test case #1557/2803" severity error;
    assert SOL = '0' report "Error in test case #1557/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1558/2803" severity error;
    assert SOR = '1' report "Error in test case #1558/2803" severity error;
    assert SOL = '0' report "Error in test case #1558/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1559/2803" severity error;
    assert SOR = '1' report "Error in test case #1559/2803" severity error;
    assert SOL = '0' report "Error in test case #1559/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1560/2803" severity error;
    assert SOR = '1' report "Error in test case #1560/2803" severity error;
    assert SOL = '0' report "Error in test case #1560/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1561/2803" severity error;
    assert SOR = '1' report "Error in test case #1561/2803" severity error;
    assert SOL = '0' report "Error in test case #1561/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1562/2803" severity error;
    assert SOR = '1' report "Error in test case #1562/2803" severity error;
    assert SOL = '0' report "Error in test case #1562/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1563/2803" severity error;
    assert SOR = '1' report "Error in test case #1563/2803" severity error;
    assert SOL = '0' report "Error in test case #1563/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1564/2803" severity error;
    assert SOR = '1' report "Error in test case #1564/2803" severity error;
    assert SOL = '0' report "Error in test case #1564/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1565/2803" severity error;
    assert SOR = '1' report "Error in test case #1565/2803" severity error;
    assert SOL = '0' report "Error in test case #1565/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1566/2803" severity error;
    assert SOR = '1' report "Error in test case #1566/2803" severity error;
    assert SOL = '0' report "Error in test case #1566/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000101" report "Error in test case #1567/2803" severity error;
    assert SOR = '1' report "Error in test case #1567/2803" severity error;
    assert SOL = '0' report "Error in test case #1567/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1568/2803" severity error;
    assert SOR = '0' report "Error in test case #1568/2803" severity error;
    assert SOL = '0' report "Error in test case #1568/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1569/2803" severity error;
    assert SOR = '0' report "Error in test case #1569/2803" severity error;
    assert SOL = '0' report "Error in test case #1569/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1570/2803" severity error;
    assert SOR = '0' report "Error in test case #1570/2803" severity error;
    assert SOL = '0' report "Error in test case #1570/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1571/2803" severity error;
    assert SOR = '0' report "Error in test case #1571/2803" severity error;
    assert SOL = '0' report "Error in test case #1571/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1572/2803" severity error;
    assert SOR = '0' report "Error in test case #1572/2803" severity error;
    assert SOL = '0' report "Error in test case #1572/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1573/2803" severity error;
    assert SOR = '0' report "Error in test case #1573/2803" severity error;
    assert SOL = '0' report "Error in test case #1573/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1574/2803" severity error;
    assert SOR = '0' report "Error in test case #1574/2803" severity error;
    assert SOL = '0' report "Error in test case #1574/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1575/2803" severity error;
    assert SOR = '0' report "Error in test case #1575/2803" severity error;
    assert SOL = '0' report "Error in test case #1575/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1576/2803" severity error;
    assert SOR = '1' report "Error in test case #1576/2803" severity error;
    assert SOL = '0' report "Error in test case #1576/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1577/2803" severity error;
    assert SOR = '1' report "Error in test case #1577/2803" severity error;
    assert SOL = '0' report "Error in test case #1577/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1578/2803" severity error;
    assert SOR = '1' report "Error in test case #1578/2803" severity error;
    assert SOL = '0' report "Error in test case #1578/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1579/2803" severity error;
    assert SOR = '1' report "Error in test case #1579/2803" severity error;
    assert SOL = '0' report "Error in test case #1579/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1580/2803" severity error;
    assert SOR = '1' report "Error in test case #1580/2803" severity error;
    assert SOL = '0' report "Error in test case #1580/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1581/2803" severity error;
    assert SOR = '1' report "Error in test case #1581/2803" severity error;
    assert SOL = '0' report "Error in test case #1581/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1582/2803" severity error;
    assert SOR = '1' report "Error in test case #1582/2803" severity error;
    assert SOL = '0' report "Error in test case #1582/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000011" report "Error in test case #1583/2803" severity error;
    assert SOR = '1' report "Error in test case #1583/2803" severity error;
    assert SOL = '0' report "Error in test case #1583/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1584/2803" severity error;
    assert SOR = '1' report "Error in test case #1584/2803" severity error;
    assert SOL = '0' report "Error in test case #1584/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1585/2803" severity error;
    assert SOR = '1' report "Error in test case #1585/2803" severity error;
    assert SOL = '0' report "Error in test case #1585/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1586/2803" severity error;
    assert SOR = '1' report "Error in test case #1586/2803" severity error;
    assert SOL = '0' report "Error in test case #1586/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1587/2803" severity error;
    assert SOR = '1' report "Error in test case #1587/2803" severity error;
    assert SOL = '0' report "Error in test case #1587/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1588/2803" severity error;
    assert SOR = '1' report "Error in test case #1588/2803" severity error;
    assert SOL = '0' report "Error in test case #1588/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1589/2803" severity error;
    assert SOR = '1' report "Error in test case #1589/2803" severity error;
    assert SOL = '0' report "Error in test case #1589/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1590/2803" severity error;
    assert SOR = '1' report "Error in test case #1590/2803" severity error;
    assert SOL = '0' report "Error in test case #1590/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1591/2803" severity error;
    assert SOR = '1' report "Error in test case #1591/2803" severity error;
    assert SOL = '0' report "Error in test case #1591/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1592/2803" severity error;
    assert SOR = '0' report "Error in test case #1592/2803" severity error;
    assert SOL = '0' report "Error in test case #1592/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1593/2803" severity error;
    assert SOR = '0' report "Error in test case #1593/2803" severity error;
    assert SOL = '0' report "Error in test case #1593/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1594/2803" severity error;
    assert SOR = '0' report "Error in test case #1594/2803" severity error;
    assert SOL = '0' report "Error in test case #1594/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1595/2803" severity error;
    assert SOR = '0' report "Error in test case #1595/2803" severity error;
    assert SOL = '0' report "Error in test case #1595/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1596/2803" severity error;
    assert SOR = '0' report "Error in test case #1596/2803" severity error;
    assert SOL = '0' report "Error in test case #1596/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1597/2803" severity error;
    assert SOR = '0' report "Error in test case #1597/2803" severity error;
    assert SOL = '0' report "Error in test case #1597/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1598/2803" severity error;
    assert SOR = '0' report "Error in test case #1598/2803" severity error;
    assert SOL = '0' report "Error in test case #1598/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000110" report "Error in test case #1599/2803" severity error;
    assert SOR = '0' report "Error in test case #1599/2803" severity error;
    assert SOL = '0' report "Error in test case #1599/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1600/2803" severity error;
    assert SOR = '1' report "Error in test case #1600/2803" severity error;
    assert SOL = '0' report "Error in test case #1600/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1601/2803" severity error;
    assert SOR = '1' report "Error in test case #1601/2803" severity error;
    assert SOL = '0' report "Error in test case #1601/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1602/2803" severity error;
    assert SOR = '1' report "Error in test case #1602/2803" severity error;
    assert SOL = '0' report "Error in test case #1602/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "011";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1603/2803" severity error;
    assert SOR = '1' report "Error in test case #1603/2803" severity error;
    assert SOL = '0' report "Error in test case #1603/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1604/2803" severity error;
    assert SOR = '1' report "Error in test case #1604/2803" severity error;
    assert SOL = '0' report "Error in test case #1604/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1605/2803" severity error;
    assert SOR = '1' report "Error in test case #1605/2803" severity error;
    assert SOL = '0' report "Error in test case #1605/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1606/2803" severity error;
    assert SOR = '1' report "Error in test case #1606/2803" severity error;
    assert SOL = '0' report "Error in test case #1606/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1607/2803" severity error;
    assert SOR = '1' report "Error in test case #1607/2803" severity error;
    assert SOL = '0' report "Error in test case #1607/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1608/2803" severity error;
    assert SOR = '1' report "Error in test case #1608/2803" severity error;
    assert SOL = '0' report "Error in test case #1608/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1609/2803" severity error;
    assert SOR = '1' report "Error in test case #1609/2803" severity error;
    assert SOL = '0' report "Error in test case #1609/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1610/2803" severity error;
    assert SOR = '1' report "Error in test case #1610/2803" severity error;
    assert SOL = '0' report "Error in test case #1610/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1611/2803" severity error;
    assert SOR = '1' report "Error in test case #1611/2803" severity error;
    assert SOL = '0' report "Error in test case #1611/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1612/2803" severity error;
    assert SOR = '1' report "Error in test case #1612/2803" severity error;
    assert SOL = '0' report "Error in test case #1612/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1613/2803" severity error;
    assert SOR = '1' report "Error in test case #1613/2803" severity error;
    assert SOL = '0' report "Error in test case #1613/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1614/2803" severity error;
    assert SOR = '1' report "Error in test case #1614/2803" severity error;
    assert SOL = '0' report "Error in test case #1614/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1615/2803" severity error;
    assert SOR = '1' report "Error in test case #1615/2803" severity error;
    assert SOL = '0' report "Error in test case #1615/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1616/2803" severity error;
    assert SOR = '1' report "Error in test case #1616/2803" severity error;
    assert SOL = '0' report "Error in test case #1616/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1617/2803" severity error;
    assert SOR = '1' report "Error in test case #1617/2803" severity error;
    assert SOL = '0' report "Error in test case #1617/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1618/2803" severity error;
    assert SOR = '1' report "Error in test case #1618/2803" severity error;
    assert SOL = '0' report "Error in test case #1618/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1619/2803" severity error;
    assert SOR = '1' report "Error in test case #1619/2803" severity error;
    assert SOL = '0' report "Error in test case #1619/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1620/2803" severity error;
    assert SOR = '1' report "Error in test case #1620/2803" severity error;
    assert SOL = '0' report "Error in test case #1620/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1621/2803" severity error;
    assert SOR = '1' report "Error in test case #1621/2803" severity error;
    assert SOL = '0' report "Error in test case #1621/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1622/2803" severity error;
    assert SOR = '1' report "Error in test case #1622/2803" severity error;
    assert SOL = '0' report "Error in test case #1622/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1623/2803" severity error;
    assert SOR = '1' report "Error in test case #1623/2803" severity error;
    assert SOL = '0' report "Error in test case #1623/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1624/2803" severity error;
    assert SOR = '1' report "Error in test case #1624/2803" severity error;
    assert SOL = '0' report "Error in test case #1624/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1625/2803" severity error;
    assert SOR = '1' report "Error in test case #1625/2803" severity error;
    assert SOL = '0' report "Error in test case #1625/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1626/2803" severity error;
    assert SOR = '1' report "Error in test case #1626/2803" severity error;
    assert SOL = '0' report "Error in test case #1626/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1627/2803" severity error;
    assert SOR = '1' report "Error in test case #1627/2803" severity error;
    assert SOL = '0' report "Error in test case #1627/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1628/2803" severity error;
    assert SOR = '1' report "Error in test case #1628/2803" severity error;
    assert SOL = '0' report "Error in test case #1628/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1629/2803" severity error;
    assert SOR = '1' report "Error in test case #1629/2803" severity error;
    assert SOL = '0' report "Error in test case #1629/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1630/2803" severity error;
    assert SOR = '1' report "Error in test case #1630/2803" severity error;
    assert SOL = '0' report "Error in test case #1630/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1631/2803" severity error;
    assert SOR = '1' report "Error in test case #1631/2803" severity error;
    assert SOL = '0' report "Error in test case #1631/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1632/2803" severity error;
    assert SOR = '1' report "Error in test case #1632/2803" severity error;
    assert SOL = '0' report "Error in test case #1632/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1633/2803" severity error;
    assert SOR = '1' report "Error in test case #1633/2803" severity error;
    assert SOL = '0' report "Error in test case #1633/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1634/2803" severity error;
    assert SOR = '1' report "Error in test case #1634/2803" severity error;
    assert SOL = '0' report "Error in test case #1634/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1635/2803" severity error;
    assert SOR = '1' report "Error in test case #1635/2803" severity error;
    assert SOL = '0' report "Error in test case #1635/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1636/2803" severity error;
    assert SOR = '1' report "Error in test case #1636/2803" severity error;
    assert SOL = '0' report "Error in test case #1636/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1637/2803" severity error;
    assert SOR = '1' report "Error in test case #1637/2803" severity error;
    assert SOL = '0' report "Error in test case #1637/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000001" report "Error in test case #1638/2803" severity error;
    assert SOR = '1' report "Error in test case #1638/2803" severity error;
    assert SOL = '0' report "Error in test case #1638/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1639/2803" severity error;
    assert SOR = '0' report "Error in test case #1639/2803" severity error;
    assert SOL = '0' report "Error in test case #1639/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1640/2803" severity error;
    assert SOR = '0' report "Error in test case #1640/2803" severity error;
    assert SOL = '0' report "Error in test case #1640/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1641/2803" severity error;
    assert SOR = '0' report "Error in test case #1641/2803" severity error;
    assert SOL = '0' report "Error in test case #1641/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1642/2803" severity error;
    assert SOR = '0' report "Error in test case #1642/2803" severity error;
    assert SOL = '0' report "Error in test case #1642/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1643/2803" severity error;
    assert SOR = '0' report "Error in test case #1643/2803" severity error;
    assert SOL = '0' report "Error in test case #1643/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1644/2803" severity error;
    assert SOR = '0' report "Error in test case #1644/2803" severity error;
    assert SOL = '0' report "Error in test case #1644/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1645/2803" severity error;
    assert SOR = '0' report "Error in test case #1645/2803" severity error;
    assert SOL = '0' report "Error in test case #1645/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1646/2803" severity error;
    assert SOR = '0' report "Error in test case #1646/2803" severity error;
    assert SOL = '0' report "Error in test case #1646/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1647/2803" severity error;
    assert SOR = '0' report "Error in test case #1647/2803" severity error;
    assert SOL = '0' report "Error in test case #1647/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1648/2803" severity error;
    assert SOR = '0' report "Error in test case #1648/2803" severity error;
    assert SOL = '0' report "Error in test case #1648/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1649/2803" severity error;
    assert SOR = '0' report "Error in test case #1649/2803" severity error;
    assert SOL = '0' report "Error in test case #1649/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1650/2803" severity error;
    assert SOR = '0' report "Error in test case #1650/2803" severity error;
    assert SOL = '0' report "Error in test case #1650/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1651/2803" severity error;
    assert SOR = '0' report "Error in test case #1651/2803" severity error;
    assert SOL = '0' report "Error in test case #1651/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1652/2803" severity error;
    assert SOR = '0' report "Error in test case #1652/2803" severity error;
    assert SOL = '0' report "Error in test case #1652/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1653/2803" severity error;
    assert SOR = '0' report "Error in test case #1653/2803" severity error;
    assert SOL = '0' report "Error in test case #1653/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1654/2803" severity error;
    assert SOR = '0' report "Error in test case #1654/2803" severity error;
    assert SOL = '0' report "Error in test case #1654/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1655/2803" severity error;
    assert SOR = '0' report "Error in test case #1655/2803" severity error;
    assert SOL = '0' report "Error in test case #1655/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1656/2803" severity error;
    assert SOR = '0' report "Error in test case #1656/2803" severity error;
    assert SOL = '0' report "Error in test case #1656/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1657/2803" severity error;
    assert SOR = '0' report "Error in test case #1657/2803" severity error;
    assert SOL = '0' report "Error in test case #1657/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1658/2803" severity error;
    assert SOR = '0' report "Error in test case #1658/2803" severity error;
    assert SOL = '0' report "Error in test case #1658/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1659/2803" severity error;
    assert SOR = '0' report "Error in test case #1659/2803" severity error;
    assert SOL = '0' report "Error in test case #1659/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1660/2803" severity error;
    assert SOR = '0' report "Error in test case #1660/2803" severity error;
    assert SOL = '0' report "Error in test case #1660/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1661/2803" severity error;
    assert SOR = '0' report "Error in test case #1661/2803" severity error;
    assert SOL = '0' report "Error in test case #1661/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1662/2803" severity error;
    assert SOR = '0' report "Error in test case #1662/2803" severity error;
    assert SOL = '0' report "Error in test case #1662/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1663/2803" severity error;
    assert SOR = '0' report "Error in test case #1663/2803" severity error;
    assert SOL = '0' report "Error in test case #1663/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1664/2803" severity error;
    assert SOR = '0' report "Error in test case #1664/2803" severity error;
    assert SOL = '0' report "Error in test case #1664/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1665/2803" severity error;
    assert SOR = '0' report "Error in test case #1665/2803" severity error;
    assert SOL = '0' report "Error in test case #1665/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1666/2803" severity error;
    assert SOR = '0' report "Error in test case #1666/2803" severity error;
    assert SOL = '0' report "Error in test case #1666/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1667/2803" severity error;
    assert SOR = '0' report "Error in test case #1667/2803" severity error;
    assert SOL = '0' report "Error in test case #1667/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1668/2803" severity error;
    assert SOR = '0' report "Error in test case #1668/2803" severity error;
    assert SOL = '0' report "Error in test case #1668/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1669/2803" severity error;
    assert SOR = '0' report "Error in test case #1669/2803" severity error;
    assert SOL = '0' report "Error in test case #1669/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1670/2803" severity error;
    assert SOR = '0' report "Error in test case #1670/2803" severity error;
    assert SOL = '0' report "Error in test case #1670/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1671/2803" severity error;
    assert SOR = '0' report "Error in test case #1671/2803" severity error;
    assert SOL = '0' report "Error in test case #1671/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1672/2803" severity error;
    assert SOR = '0' report "Error in test case #1672/2803" severity error;
    assert SOL = '0' report "Error in test case #1672/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1673/2803" severity error;
    assert SOR = '0' report "Error in test case #1673/2803" severity error;
    assert SOL = '0' report "Error in test case #1673/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1674/2803" severity error;
    assert SOR = '0' report "Error in test case #1674/2803" severity error;
    assert SOL = '0' report "Error in test case #1674/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1675/2803" severity error;
    assert SOR = '0' report "Error in test case #1675/2803" severity error;
    assert SOL = '0' report "Error in test case #1675/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1676/2803" severity error;
    assert SOR = '0' report "Error in test case #1676/2803" severity error;
    assert SOL = '0' report "Error in test case #1676/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1677/2803" severity error;
    assert SOR = '0' report "Error in test case #1677/2803" severity error;
    assert SOL = '0' report "Error in test case #1677/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1678/2803" severity error;
    assert SOR = '0' report "Error in test case #1678/2803" severity error;
    assert SOL = '0' report "Error in test case #1678/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1679/2803" severity error;
    assert SOR = '0' report "Error in test case #1679/2803" severity error;
    assert SOL = '0' report "Error in test case #1679/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1680/2803" severity error;
    assert SOR = '0' report "Error in test case #1680/2803" severity error;
    assert SOL = '0' report "Error in test case #1680/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1681/2803" severity error;
    assert SOR = '0' report "Error in test case #1681/2803" severity error;
    assert SOL = '0' report "Error in test case #1681/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1682/2803" severity error;
    assert SOR = '0' report "Error in test case #1682/2803" severity error;
    assert SOL = '0' report "Error in test case #1682/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1683/2803" severity error;
    assert SOR = '0' report "Error in test case #1683/2803" severity error;
    assert SOL = '0' report "Error in test case #1683/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1684/2803" severity error;
    assert SOR = '0' report "Error in test case #1684/2803" severity error;
    assert SOL = '0' report "Error in test case #1684/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1685/2803" severity error;
    assert SOR = '0' report "Error in test case #1685/2803" severity error;
    assert SOL = '0' report "Error in test case #1685/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1686/2803" severity error;
    assert SOR = '0' report "Error in test case #1686/2803" severity error;
    assert SOL = '0' report "Error in test case #1686/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1687/2803" severity error;
    assert SOR = '0' report "Error in test case #1687/2803" severity error;
    assert SOL = '0' report "Error in test case #1687/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1688/2803" severity error;
    assert SOR = '0' report "Error in test case #1688/2803" severity error;
    assert SOL = '0' report "Error in test case #1688/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1689/2803" severity error;
    assert SOR = '0' report "Error in test case #1689/2803" severity error;
    assert SOL = '0' report "Error in test case #1689/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1690/2803" severity error;
    assert SOR = '0' report "Error in test case #1690/2803" severity error;
    assert SOL = '0' report "Error in test case #1690/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1691/2803" severity error;
    assert SOR = '0' report "Error in test case #1691/2803" severity error;
    assert SOL = '0' report "Error in test case #1691/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1692/2803" severity error;
    assert SOR = '0' report "Error in test case #1692/2803" severity error;
    assert SOL = '0' report "Error in test case #1692/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1693/2803" severity error;
    assert SOR = '0' report "Error in test case #1693/2803" severity error;
    assert SOL = '0' report "Error in test case #1693/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1694/2803" severity error;
    assert SOR = '0' report "Error in test case #1694/2803" severity error;
    assert SOL = '0' report "Error in test case #1694/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1695/2803" severity error;
    assert SOR = '0' report "Error in test case #1695/2803" severity error;
    assert SOL = '0' report "Error in test case #1695/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1696/2803" severity error;
    assert SOR = '0' report "Error in test case #1696/2803" severity error;
    assert SOL = '0' report "Error in test case #1696/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1697/2803" severity error;
    assert SOR = '0' report "Error in test case #1697/2803" severity error;
    assert SOL = '0' report "Error in test case #1697/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1698/2803" severity error;
    assert SOR = '0' report "Error in test case #1698/2803" severity error;
    assert SOL = '0' report "Error in test case #1698/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1699/2803" severity error;
    assert SOR = '0' report "Error in test case #1699/2803" severity error;
    assert SOL = '0' report "Error in test case #1699/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1700/2803" severity error;
    assert SOR = '0' report "Error in test case #1700/2803" severity error;
    assert SOL = '0' report "Error in test case #1700/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1701/2803" severity error;
    assert SOR = '0' report "Error in test case #1701/2803" severity error;
    assert SOL = '0' report "Error in test case #1701/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1702/2803" severity error;
    assert SOR = '0' report "Error in test case #1702/2803" severity error;
    assert SOL = '0' report "Error in test case #1702/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1703/2803" severity error;
    assert SOR = '0' report "Error in test case #1703/2803" severity error;
    assert SOL = '0' report "Error in test case #1703/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1704/2803" severity error;
    assert SOR = '0' report "Error in test case #1704/2803" severity error;
    assert SOL = '0' report "Error in test case #1704/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1705/2803" severity error;
    assert SOR = '0' report "Error in test case #1705/2803" severity error;
    assert SOL = '0' report "Error in test case #1705/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1706/2803" severity error;
    assert SOR = '0' report "Error in test case #1706/2803" severity error;
    assert SOL = '0' report "Error in test case #1706/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1707/2803" severity error;
    assert SOR = '0' report "Error in test case #1707/2803" severity error;
    assert SOL = '0' report "Error in test case #1707/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1708/2803" severity error;
    assert SOR = '0' report "Error in test case #1708/2803" severity error;
    assert SOL = '0' report "Error in test case #1708/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1709/2803" severity error;
    assert SOR = '0' report "Error in test case #1709/2803" severity error;
    assert SOL = '0' report "Error in test case #1709/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1710/2803" severity error;
    assert SOR = '0' report "Error in test case #1710/2803" severity error;
    assert SOL = '0' report "Error in test case #1710/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1711/2803" severity error;
    assert SOR = '0' report "Error in test case #1711/2803" severity error;
    assert SOL = '0' report "Error in test case #1711/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1712/2803" severity error;
    assert SOR = '0' report "Error in test case #1712/2803" severity error;
    assert SOL = '0' report "Error in test case #1712/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1713/2803" severity error;
    assert SOR = '0' report "Error in test case #1713/2803" severity error;
    assert SOL = '0' report "Error in test case #1713/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1714/2803" severity error;
    assert SOR = '0' report "Error in test case #1714/2803" severity error;
    assert SOL = '0' report "Error in test case #1714/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1715/2803" severity error;
    assert SOR = '0' report "Error in test case #1715/2803" severity error;
    assert SOL = '0' report "Error in test case #1715/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1716/2803" severity error;
    assert SOR = '0' report "Error in test case #1716/2803" severity error;
    assert SOL = '0' report "Error in test case #1716/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1717/2803" severity error;
    assert SOR = '0' report "Error in test case #1717/2803" severity error;
    assert SOL = '0' report "Error in test case #1717/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1718/2803" severity error;
    assert SOR = '0' report "Error in test case #1718/2803" severity error;
    assert SOL = '0' report "Error in test case #1718/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1719/2803" severity error;
    assert SOR = '0' report "Error in test case #1719/2803" severity error;
    assert SOL = '0' report "Error in test case #1719/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1720/2803" severity error;
    assert SOR = '0' report "Error in test case #1720/2803" severity error;
    assert SOL = '0' report "Error in test case #1720/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1721/2803" severity error;
    assert SOR = '0' report "Error in test case #1721/2803" severity error;
    assert SOL = '0' report "Error in test case #1721/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1722/2803" severity error;
    assert SOR = '0' report "Error in test case #1722/2803" severity error;
    assert SOL = '0' report "Error in test case #1722/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1723/2803" severity error;
    assert SOR = '0' report "Error in test case #1723/2803" severity error;
    assert SOL = '0' report "Error in test case #1723/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1724/2803" severity error;
    assert SOR = '0' report "Error in test case #1724/2803" severity error;
    assert SOL = '0' report "Error in test case #1724/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1725/2803" severity error;
    assert SOR = '0' report "Error in test case #1725/2803" severity error;
    assert SOL = '0' report "Error in test case #1725/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1726/2803" severity error;
    assert SOR = '0' report "Error in test case #1726/2803" severity error;
    assert SOL = '0' report "Error in test case #1726/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1727/2803" severity error;
    assert SOR = '1' report "Error in test case #1727/2803" severity error;
    assert SOL = '1' report "Error in test case #1727/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1728/2803" severity error;
    assert SOR = '1' report "Error in test case #1728/2803" severity error;
    assert SOL = '1' report "Error in test case #1728/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1729/2803" severity error;
    assert SOR = '1' report "Error in test case #1729/2803" severity error;
    assert SOL = '1' report "Error in test case #1729/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1730/2803" severity error;
    assert SOR = '1' report "Error in test case #1730/2803" severity error;
    assert SOL = '1' report "Error in test case #1730/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1731/2803" severity error;
    assert SOR = '1' report "Error in test case #1731/2803" severity error;
    assert SOL = '1' report "Error in test case #1731/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1732/2803" severity error;
    assert SOR = '1' report "Error in test case #1732/2803" severity error;
    assert SOL = '1' report "Error in test case #1732/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1733/2803" severity error;
    assert SOR = '1' report "Error in test case #1733/2803" severity error;
    assert SOL = '1' report "Error in test case #1733/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1734/2803" severity error;
    assert SOR = '1' report "Error in test case #1734/2803" severity error;
    assert SOL = '1' report "Error in test case #1734/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1735/2803" severity error;
    assert SOR = '1' report "Error in test case #1735/2803" severity error;
    assert SOL = '1' report "Error in test case #1735/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1736/2803" severity error;
    assert SOR = '1' report "Error in test case #1736/2803" severity error;
    assert SOL = '1' report "Error in test case #1736/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1737/2803" severity error;
    assert SOR = '1' report "Error in test case #1737/2803" severity error;
    assert SOL = '1' report "Error in test case #1737/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1738/2803" severity error;
    assert SOR = '1' report "Error in test case #1738/2803" severity error;
    assert SOL = '1' report "Error in test case #1738/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1739/2803" severity error;
    assert SOR = '1' report "Error in test case #1739/2803" severity error;
    assert SOL = '1' report "Error in test case #1739/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1740/2803" severity error;
    assert SOR = '1' report "Error in test case #1740/2803" severity error;
    assert SOL = '1' report "Error in test case #1740/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1741/2803" severity error;
    assert SOR = '1' report "Error in test case #1741/2803" severity error;
    assert SOL = '1' report "Error in test case #1741/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1742/2803" severity error;
    assert SOR = '1' report "Error in test case #1742/2803" severity error;
    assert SOL = '1' report "Error in test case #1742/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1743/2803" severity error;
    assert SOR = '1' report "Error in test case #1743/2803" severity error;
    assert SOL = '1' report "Error in test case #1743/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1744/2803" severity error;
    assert SOR = '1' report "Error in test case #1744/2803" severity error;
    assert SOL = '1' report "Error in test case #1744/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1745/2803" severity error;
    assert SOR = '1' report "Error in test case #1745/2803" severity error;
    assert SOL = '1' report "Error in test case #1745/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1746/2803" severity error;
    assert SOR = '1' report "Error in test case #1746/2803" severity error;
    assert SOL = '1' report "Error in test case #1746/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1747/2803" severity error;
    assert SOR = '1' report "Error in test case #1747/2803" severity error;
    assert SOL = '1' report "Error in test case #1747/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1748/2803" severity error;
    assert SOR = '1' report "Error in test case #1748/2803" severity error;
    assert SOL = '1' report "Error in test case #1748/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1749/2803" severity error;
    assert SOR = '1' report "Error in test case #1749/2803" severity error;
    assert SOL = '1' report "Error in test case #1749/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1750/2803" severity error;
    assert SOR = '1' report "Error in test case #1750/2803" severity error;
    assert SOL = '1' report "Error in test case #1750/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1751/2803" severity error;
    assert SOR = '1' report "Error in test case #1751/2803" severity error;
    assert SOL = '1' report "Error in test case #1751/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1752/2803" severity error;
    assert SOR = '1' report "Error in test case #1752/2803" severity error;
    assert SOL = '1' report "Error in test case #1752/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1753/2803" severity error;
    assert SOR = '1' report "Error in test case #1753/2803" severity error;
    assert SOL = '1' report "Error in test case #1753/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1754/2803" severity error;
    assert SOR = '1' report "Error in test case #1754/2803" severity error;
    assert SOL = '1' report "Error in test case #1754/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1755/2803" severity error;
    assert SOR = '1' report "Error in test case #1755/2803" severity error;
    assert SOL = '1' report "Error in test case #1755/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1756/2803" severity error;
    assert SOR = '1' report "Error in test case #1756/2803" severity error;
    assert SOL = '1' report "Error in test case #1756/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1757/2803" severity error;
    assert SOR = '1' report "Error in test case #1757/2803" severity error;
    assert SOL = '1' report "Error in test case #1757/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1758/2803" severity error;
    assert SOR = '1' report "Error in test case #1758/2803" severity error;
    assert SOL = '1' report "Error in test case #1758/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1759/2803" severity error;
    assert SOR = '1' report "Error in test case #1759/2803" severity error;
    assert SOL = '1' report "Error in test case #1759/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1760/2803" severity error;
    assert SOR = '1' report "Error in test case #1760/2803" severity error;
    assert SOL = '1' report "Error in test case #1760/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1761/2803" severity error;
    assert SOR = '1' report "Error in test case #1761/2803" severity error;
    assert SOL = '1' report "Error in test case #1761/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1762/2803" severity error;
    assert SOR = '1' report "Error in test case #1762/2803" severity error;
    assert SOL = '1' report "Error in test case #1762/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1763/2803" severity error;
    assert SOR = '1' report "Error in test case #1763/2803" severity error;
    assert SOL = '1' report "Error in test case #1763/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1764/2803" severity error;
    assert SOR = '1' report "Error in test case #1764/2803" severity error;
    assert SOL = '1' report "Error in test case #1764/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1765/2803" severity error;
    assert SOR = '1' report "Error in test case #1765/2803" severity error;
    assert SOL = '1' report "Error in test case #1765/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1766/2803" severity error;
    assert SOR = '1' report "Error in test case #1766/2803" severity error;
    assert SOL = '1' report "Error in test case #1766/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1767/2803" severity error;
    assert SOR = '1' report "Error in test case #1767/2803" severity error;
    assert SOL = '1' report "Error in test case #1767/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1768/2803" severity error;
    assert SOR = '1' report "Error in test case #1768/2803" severity error;
    assert SOL = '1' report "Error in test case #1768/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1769/2803" severity error;
    assert SOR = '1' report "Error in test case #1769/2803" severity error;
    assert SOL = '1' report "Error in test case #1769/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1770/2803" severity error;
    assert SOR = '1' report "Error in test case #1770/2803" severity error;
    assert SOL = '1' report "Error in test case #1770/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1771/2803" severity error;
    assert SOR = '1' report "Error in test case #1771/2803" severity error;
    assert SOL = '1' report "Error in test case #1771/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1772/2803" severity error;
    assert SOR = '1' report "Error in test case #1772/2803" severity error;
    assert SOL = '1' report "Error in test case #1772/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1773/2803" severity error;
    assert SOR = '1' report "Error in test case #1773/2803" severity error;
    assert SOL = '1' report "Error in test case #1773/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1774/2803" severity error;
    assert SOR = '1' report "Error in test case #1774/2803" severity error;
    assert SOL = '1' report "Error in test case #1774/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1775/2803" severity error;
    assert SOR = '1' report "Error in test case #1775/2803" severity error;
    assert SOL = '1' report "Error in test case #1775/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1776/2803" severity error;
    assert SOR = '1' report "Error in test case #1776/2803" severity error;
    assert SOL = '1' report "Error in test case #1776/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1777/2803" severity error;
    assert SOR = '1' report "Error in test case #1777/2803" severity error;
    assert SOL = '1' report "Error in test case #1777/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1778/2803" severity error;
    assert SOR = '1' report "Error in test case #1778/2803" severity error;
    assert SOL = '1' report "Error in test case #1778/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1779/2803" severity error;
    assert SOR = '1' report "Error in test case #1779/2803" severity error;
    assert SOL = '1' report "Error in test case #1779/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1780/2803" severity error;
    assert SOR = '1' report "Error in test case #1780/2803" severity error;
    assert SOL = '1' report "Error in test case #1780/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1781/2803" severity error;
    assert SOR = '1' report "Error in test case #1781/2803" severity error;
    assert SOL = '1' report "Error in test case #1781/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1782/2803" severity error;
    assert SOR = '1' report "Error in test case #1782/2803" severity error;
    assert SOL = '1' report "Error in test case #1782/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1783/2803" severity error;
    assert SOR = '1' report "Error in test case #1783/2803" severity error;
    assert SOL = '1' report "Error in test case #1783/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1784/2803" severity error;
    assert SOR = '1' report "Error in test case #1784/2803" severity error;
    assert SOL = '1' report "Error in test case #1784/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1785/2803" severity error;
    assert SOR = '1' report "Error in test case #1785/2803" severity error;
    assert SOL = '1' report "Error in test case #1785/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1786/2803" severity error;
    assert SOR = '1' report "Error in test case #1786/2803" severity error;
    assert SOL = '1' report "Error in test case #1786/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1787/2803" severity error;
    assert SOR = '1' report "Error in test case #1787/2803" severity error;
    assert SOL = '1' report "Error in test case #1787/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1788/2803" severity error;
    assert SOR = '1' report "Error in test case #1788/2803" severity error;
    assert SOL = '1' report "Error in test case #1788/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1789/2803" severity error;
    assert SOR = '1' report "Error in test case #1789/2803" severity error;
    assert SOL = '1' report "Error in test case #1789/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1790/2803" severity error;
    assert SOR = '1' report "Error in test case #1790/2803" severity error;
    assert SOL = '1' report "Error in test case #1790/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1791/2803" severity error;
    assert SOR = '1' report "Error in test case #1791/2803" severity error;
    assert SOL = '1' report "Error in test case #1791/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1792/2803" severity error;
    assert SOR = '1' report "Error in test case #1792/2803" severity error;
    assert SOL = '1' report "Error in test case #1792/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1793/2803" severity error;
    assert SOR = '1' report "Error in test case #1793/2803" severity error;
    assert SOL = '1' report "Error in test case #1793/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1794/2803" severity error;
    assert SOR = '1' report "Error in test case #1794/2803" severity error;
    assert SOL = '1' report "Error in test case #1794/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1795/2803" severity error;
    assert SOR = '1' report "Error in test case #1795/2803" severity error;
    assert SOL = '1' report "Error in test case #1795/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1796/2803" severity error;
    assert SOR = '1' report "Error in test case #1796/2803" severity error;
    assert SOL = '1' report "Error in test case #1796/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1797/2803" severity error;
    assert SOR = '1' report "Error in test case #1797/2803" severity error;
    assert SOL = '1' report "Error in test case #1797/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1798/2803" severity error;
    assert SOR = '1' report "Error in test case #1798/2803" severity error;
    assert SOL = '1' report "Error in test case #1798/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1799/2803" severity error;
    assert SOR = '1' report "Error in test case #1799/2803" severity error;
    assert SOL = '1' report "Error in test case #1799/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1800/2803" severity error;
    assert SOR = '1' report "Error in test case #1800/2803" severity error;
    assert SOL = '1' report "Error in test case #1800/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1801/2803" severity error;
    assert SOR = '1' report "Error in test case #1801/2803" severity error;
    assert SOL = '1' report "Error in test case #1801/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1802/2803" severity error;
    assert SOR = '1' report "Error in test case #1802/2803" severity error;
    assert SOL = '1' report "Error in test case #1802/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1803/2803" severity error;
    assert SOR = '1' report "Error in test case #1803/2803" severity error;
    assert SOL = '1' report "Error in test case #1803/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1804/2803" severity error;
    assert SOR = '1' report "Error in test case #1804/2803" severity error;
    assert SOL = '1' report "Error in test case #1804/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1805/2803" severity error;
    assert SOR = '1' report "Error in test case #1805/2803" severity error;
    assert SOL = '1' report "Error in test case #1805/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1806/2803" severity error;
    assert SOR = '1' report "Error in test case #1806/2803" severity error;
    assert SOL = '1' report "Error in test case #1806/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1807/2803" severity error;
    assert SOR = '1' report "Error in test case #1807/2803" severity error;
    assert SOL = '1' report "Error in test case #1807/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1808/2803" severity error;
    assert SOR = '1' report "Error in test case #1808/2803" severity error;
    assert SOL = '1' report "Error in test case #1808/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1809/2803" severity error;
    assert SOR = '1' report "Error in test case #1809/2803" severity error;
    assert SOL = '1' report "Error in test case #1809/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1810/2803" severity error;
    assert SOR = '1' report "Error in test case #1810/2803" severity error;
    assert SOL = '1' report "Error in test case #1810/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1811/2803" severity error;
    assert SOR = '1' report "Error in test case #1811/2803" severity error;
    assert SOL = '1' report "Error in test case #1811/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1812/2803" severity error;
    assert SOR = '1' report "Error in test case #1812/2803" severity error;
    assert SOL = '1' report "Error in test case #1812/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1813/2803" severity error;
    assert SOR = '1' report "Error in test case #1813/2803" severity error;
    assert SOL = '1' report "Error in test case #1813/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1814/2803" severity error;
    assert SOR = '1' report "Error in test case #1814/2803" severity error;
    assert SOL = '1' report "Error in test case #1814/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1815/2803" severity error;
    assert SOR = '1' report "Error in test case #1815/2803" severity error;
    assert SOL = '1' report "Error in test case #1815/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1816/2803" severity error;
    assert SOR = '1' report "Error in test case #1816/2803" severity error;
    assert SOL = '1' report "Error in test case #1816/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1817/2803" severity error;
    assert SOR = '1' report "Error in test case #1817/2803" severity error;
    assert SOL = '1' report "Error in test case #1817/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1818/2803" severity error;
    assert SOR = '1' report "Error in test case #1818/2803" severity error;
    assert SOL = '1' report "Error in test case #1818/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1819/2803" severity error;
    assert SOR = '1' report "Error in test case #1819/2803" severity error;
    assert SOL = '1' report "Error in test case #1819/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1820/2803" severity error;
    assert SOR = '1' report "Error in test case #1820/2803" severity error;
    assert SOL = '1' report "Error in test case #1820/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1821/2803" severity error;
    assert SOR = '1' report "Error in test case #1821/2803" severity error;
    assert SOL = '1' report "Error in test case #1821/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1822/2803" severity error;
    assert SOR = '1' report "Error in test case #1822/2803" severity error;
    assert SOL = '1' report "Error in test case #1822/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1823/2803" severity error;
    assert SOR = '1' report "Error in test case #1823/2803" severity error;
    assert SOL = '1' report "Error in test case #1823/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1824/2803" severity error;
    assert SOR = '1' report "Error in test case #1824/2803" severity error;
    assert SOL = '1' report "Error in test case #1824/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1825/2803" severity error;
    assert SOR = '1' report "Error in test case #1825/2803" severity error;
    assert SOL = '1' report "Error in test case #1825/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1826/2803" severity error;
    assert SOR = '1' report "Error in test case #1826/2803" severity error;
    assert SOL = '1' report "Error in test case #1826/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1827/2803" severity error;
    assert SOR = '1' report "Error in test case #1827/2803" severity error;
    assert SOL = '1' report "Error in test case #1827/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1828/2803" severity error;
    assert SOR = '1' report "Error in test case #1828/2803" severity error;
    assert SOL = '1' report "Error in test case #1828/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1829/2803" severity error;
    assert SOR = '1' report "Error in test case #1829/2803" severity error;
    assert SOL = '1' report "Error in test case #1829/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1830/2803" severity error;
    assert SOR = '1' report "Error in test case #1830/2803" severity error;
    assert SOL = '1' report "Error in test case #1830/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1831/2803" severity error;
    assert SOR = '1' report "Error in test case #1831/2803" severity error;
    assert SOL = '1' report "Error in test case #1831/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1832/2803" severity error;
    assert SOR = '1' report "Error in test case #1832/2803" severity error;
    assert SOL = '1' report "Error in test case #1832/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1833/2803" severity error;
    assert SOR = '1' report "Error in test case #1833/2803" severity error;
    assert SOL = '1' report "Error in test case #1833/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1834/2803" severity error;
    assert SOR = '1' report "Error in test case #1834/2803" severity error;
    assert SOL = '1' report "Error in test case #1834/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1835/2803" severity error;
    assert SOR = '1' report "Error in test case #1835/2803" severity error;
    assert SOL = '1' report "Error in test case #1835/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1836/2803" severity error;
    assert SOR = '1' report "Error in test case #1836/2803" severity error;
    assert SOL = '1' report "Error in test case #1836/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1837/2803" severity error;
    assert SOR = '1' report "Error in test case #1837/2803" severity error;
    assert SOL = '1' report "Error in test case #1837/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1838/2803" severity error;
    assert SOR = '1' report "Error in test case #1838/2803" severity error;
    assert SOL = '1' report "Error in test case #1838/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1839/2803" severity error;
    assert SOR = '1' report "Error in test case #1839/2803" severity error;
    assert SOL = '1' report "Error in test case #1839/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1840/2803" severity error;
    assert SOR = '1' report "Error in test case #1840/2803" severity error;
    assert SOL = '1' report "Error in test case #1840/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1841/2803" severity error;
    assert SOR = '1' report "Error in test case #1841/2803" severity error;
    assert SOL = '1' report "Error in test case #1841/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1842/2803" severity error;
    assert SOR = '1' report "Error in test case #1842/2803" severity error;
    assert SOL = '1' report "Error in test case #1842/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1843/2803" severity error;
    assert SOR = '1' report "Error in test case #1843/2803" severity error;
    assert SOL = '1' report "Error in test case #1843/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1844/2803" severity error;
    assert SOR = '1' report "Error in test case #1844/2803" severity error;
    assert SOL = '1' report "Error in test case #1844/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1845/2803" severity error;
    assert SOR = '1' report "Error in test case #1845/2803" severity error;
    assert SOL = '1' report "Error in test case #1845/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1846/2803" severity error;
    assert SOR = '1' report "Error in test case #1846/2803" severity error;
    assert SOL = '1' report "Error in test case #1846/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1847/2803" severity error;
    assert SOR = '1' report "Error in test case #1847/2803" severity error;
    assert SOL = '1' report "Error in test case #1847/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1848/2803" severity error;
    assert SOR = '1' report "Error in test case #1848/2803" severity error;
    assert SOL = '1' report "Error in test case #1848/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1849/2803" severity error;
    assert SOR = '1' report "Error in test case #1849/2803" severity error;
    assert SOL = '1' report "Error in test case #1849/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1850/2803" severity error;
    assert SOR = '1' report "Error in test case #1850/2803" severity error;
    assert SOL = '1' report "Error in test case #1850/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1851/2803" severity error;
    assert SOR = '1' report "Error in test case #1851/2803" severity error;
    assert SOL = '1' report "Error in test case #1851/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1852/2803" severity error;
    assert SOR = '1' report "Error in test case #1852/2803" severity error;
    assert SOL = '1' report "Error in test case #1852/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1853/2803" severity error;
    assert SOR = '1' report "Error in test case #1853/2803" severity error;
    assert SOL = '1' report "Error in test case #1853/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1854/2803" severity error;
    assert SOR = '1' report "Error in test case #1854/2803" severity error;
    assert SOL = '1' report "Error in test case #1854/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1855/2803" severity error;
    assert SOR = '1' report "Error in test case #1855/2803" severity error;
    assert SOL = '1' report "Error in test case #1855/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1856/2803" severity error;
    assert SOR = '1' report "Error in test case #1856/2803" severity error;
    assert SOL = '1' report "Error in test case #1856/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1857/2803" severity error;
    assert SOR = '1' report "Error in test case #1857/2803" severity error;
    assert SOL = '1' report "Error in test case #1857/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1858/2803" severity error;
    assert SOR = '1' report "Error in test case #1858/2803" severity error;
    assert SOL = '1' report "Error in test case #1858/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1859/2803" severity error;
    assert SOR = '1' report "Error in test case #1859/2803" severity error;
    assert SOL = '1' report "Error in test case #1859/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1860/2803" severity error;
    assert SOR = '1' report "Error in test case #1860/2803" severity error;
    assert SOL = '1' report "Error in test case #1860/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1861/2803" severity error;
    assert SOR = '1' report "Error in test case #1861/2803" severity error;
    assert SOL = '1' report "Error in test case #1861/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1862/2803" severity error;
    assert SOR = '1' report "Error in test case #1862/2803" severity error;
    assert SOL = '1' report "Error in test case #1862/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1863/2803" severity error;
    assert SOR = '1' report "Error in test case #1863/2803" severity error;
    assert SOL = '1' report "Error in test case #1863/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1864/2803" severity error;
    assert SOR = '1' report "Error in test case #1864/2803" severity error;
    assert SOL = '1' report "Error in test case #1864/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1865/2803" severity error;
    assert SOR = '1' report "Error in test case #1865/2803" severity error;
    assert SOL = '1' report "Error in test case #1865/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1866/2803" severity error;
    assert SOR = '1' report "Error in test case #1866/2803" severity error;
    assert SOL = '1' report "Error in test case #1866/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1867/2803" severity error;
    assert SOR = '1' report "Error in test case #1867/2803" severity error;
    assert SOL = '1' report "Error in test case #1867/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1868/2803" severity error;
    assert SOR = '1' report "Error in test case #1868/2803" severity error;
    assert SOL = '1' report "Error in test case #1868/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1869/2803" severity error;
    assert SOR = '1' report "Error in test case #1869/2803" severity error;
    assert SOL = '1' report "Error in test case #1869/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1870/2803" severity error;
    assert SOR = '1' report "Error in test case #1870/2803" severity error;
    assert SOL = '1' report "Error in test case #1870/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1871/2803" severity error;
    assert SOR = '1' report "Error in test case #1871/2803" severity error;
    assert SOL = '1' report "Error in test case #1871/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1872/2803" severity error;
    assert SOR = '1' report "Error in test case #1872/2803" severity error;
    assert SOL = '1' report "Error in test case #1872/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1873/2803" severity error;
    assert SOR = '1' report "Error in test case #1873/2803" severity error;
    assert SOL = '1' report "Error in test case #1873/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1874/2803" severity error;
    assert SOR = '1' report "Error in test case #1874/2803" severity error;
    assert SOL = '1' report "Error in test case #1874/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1875/2803" severity error;
    assert SOR = '1' report "Error in test case #1875/2803" severity error;
    assert SOL = '1' report "Error in test case #1875/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1876/2803" severity error;
    assert SOR = '1' report "Error in test case #1876/2803" severity error;
    assert SOL = '1' report "Error in test case #1876/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1877/2803" severity error;
    assert SOR = '1' report "Error in test case #1877/2803" severity error;
    assert SOL = '1' report "Error in test case #1877/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1878/2803" severity error;
    assert SOR = '1' report "Error in test case #1878/2803" severity error;
    assert SOL = '1' report "Error in test case #1878/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1879/2803" severity error;
    assert SOR = '1' report "Error in test case #1879/2803" severity error;
    assert SOL = '1' report "Error in test case #1879/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1880/2803" severity error;
    assert SOR = '1' report "Error in test case #1880/2803" severity error;
    assert SOL = '1' report "Error in test case #1880/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1881/2803" severity error;
    assert SOR = '1' report "Error in test case #1881/2803" severity error;
    assert SOL = '1' report "Error in test case #1881/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1882/2803" severity error;
    assert SOR = '1' report "Error in test case #1882/2803" severity error;
    assert SOL = '1' report "Error in test case #1882/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1883/2803" severity error;
    assert SOR = '1' report "Error in test case #1883/2803" severity error;
    assert SOL = '1' report "Error in test case #1883/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1884/2803" severity error;
    assert SOR = '1' report "Error in test case #1884/2803" severity error;
    assert SOL = '1' report "Error in test case #1884/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1885/2803" severity error;
    assert SOR = '1' report "Error in test case #1885/2803" severity error;
    assert SOL = '1' report "Error in test case #1885/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1886/2803" severity error;
    assert SOR = '1' report "Error in test case #1886/2803" severity error;
    assert SOL = '1' report "Error in test case #1886/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1887/2803" severity error;
    assert SOR = '1' report "Error in test case #1887/2803" severity error;
    assert SOL = '1' report "Error in test case #1887/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1888/2803" severity error;
    assert SOR = '1' report "Error in test case #1888/2803" severity error;
    assert SOL = '1' report "Error in test case #1888/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1889/2803" severity error;
    assert SOR = '1' report "Error in test case #1889/2803" severity error;
    assert SOL = '1' report "Error in test case #1889/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1890/2803" severity error;
    assert SOR = '1' report "Error in test case #1890/2803" severity error;
    assert SOL = '1' report "Error in test case #1890/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1891/2803" severity error;
    assert SOR = '1' report "Error in test case #1891/2803" severity error;
    assert SOL = '1' report "Error in test case #1891/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1892/2803" severity error;
    assert SOR = '1' report "Error in test case #1892/2803" severity error;
    assert SOL = '1' report "Error in test case #1892/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1893/2803" severity error;
    assert SOR = '1' report "Error in test case #1893/2803" severity error;
    assert SOL = '1' report "Error in test case #1893/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1894/2803" severity error;
    assert SOR = '1' report "Error in test case #1894/2803" severity error;
    assert SOL = '1' report "Error in test case #1894/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1895/2803" severity error;
    assert SOR = '1' report "Error in test case #1895/2803" severity error;
    assert SOL = '1' report "Error in test case #1895/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1896/2803" severity error;
    assert SOR = '1' report "Error in test case #1896/2803" severity error;
    assert SOL = '1' report "Error in test case #1896/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1897/2803" severity error;
    assert SOR = '1' report "Error in test case #1897/2803" severity error;
    assert SOL = '1' report "Error in test case #1897/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1898/2803" severity error;
    assert SOR = '1' report "Error in test case #1898/2803" severity error;
    assert SOL = '1' report "Error in test case #1898/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1899/2803" severity error;
    assert SOR = '1' report "Error in test case #1899/2803" severity error;
    assert SOL = '1' report "Error in test case #1899/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1900/2803" severity error;
    assert SOR = '1' report "Error in test case #1900/2803" severity error;
    assert SOL = '1' report "Error in test case #1900/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1901/2803" severity error;
    assert SOR = '1' report "Error in test case #1901/2803" severity error;
    assert SOL = '1' report "Error in test case #1901/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1902/2803" severity error;
    assert SOR = '1' report "Error in test case #1902/2803" severity error;
    assert SOL = '1' report "Error in test case #1902/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1903/2803" severity error;
    assert SOR = '1' report "Error in test case #1903/2803" severity error;
    assert SOL = '1' report "Error in test case #1903/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1904/2803" severity error;
    assert SOR = '1' report "Error in test case #1904/2803" severity error;
    assert SOL = '1' report "Error in test case #1904/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1905/2803" severity error;
    assert SOR = '1' report "Error in test case #1905/2803" severity error;
    assert SOL = '1' report "Error in test case #1905/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1906/2803" severity error;
    assert SOR = '1' report "Error in test case #1906/2803" severity error;
    assert SOL = '1' report "Error in test case #1906/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1907/2803" severity error;
    assert SOR = '1' report "Error in test case #1907/2803" severity error;
    assert SOL = '1' report "Error in test case #1907/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1908/2803" severity error;
    assert SOR = '1' report "Error in test case #1908/2803" severity error;
    assert SOL = '1' report "Error in test case #1908/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1909/2803" severity error;
    assert SOR = '1' report "Error in test case #1909/2803" severity error;
    assert SOL = '1' report "Error in test case #1909/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1910/2803" severity error;
    assert SOR = '1' report "Error in test case #1910/2803" severity error;
    assert SOL = '1' report "Error in test case #1910/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1911/2803" severity error;
    assert SOR = '1' report "Error in test case #1911/2803" severity error;
    assert SOL = '1' report "Error in test case #1911/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1912/2803" severity error;
    assert SOR = '1' report "Error in test case #1912/2803" severity error;
    assert SOL = '1' report "Error in test case #1912/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1913/2803" severity error;
    assert SOR = '1' report "Error in test case #1913/2803" severity error;
    assert SOL = '1' report "Error in test case #1913/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1914/2803" severity error;
    assert SOR = '1' report "Error in test case #1914/2803" severity error;
    assert SOL = '1' report "Error in test case #1914/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1915/2803" severity error;
    assert SOR = '1' report "Error in test case #1915/2803" severity error;
    assert SOL = '1' report "Error in test case #1915/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1916/2803" severity error;
    assert SOR = '1' report "Error in test case #1916/2803" severity error;
    assert SOL = '1' report "Error in test case #1916/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1917/2803" severity error;
    assert SOR = '1' report "Error in test case #1917/2803" severity error;
    assert SOL = '1' report "Error in test case #1917/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1918/2803" severity error;
    assert SOR = '1' report "Error in test case #1918/2803" severity error;
    assert SOL = '1' report "Error in test case #1918/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1919/2803" severity error;
    assert SOR = '1' report "Error in test case #1919/2803" severity error;
    assert SOL = '1' report "Error in test case #1919/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1920/2803" severity error;
    assert SOR = '1' report "Error in test case #1920/2803" severity error;
    assert SOL = '1' report "Error in test case #1920/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1921/2803" severity error;
    assert SOR = '1' report "Error in test case #1921/2803" severity error;
    assert SOL = '1' report "Error in test case #1921/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1922/2803" severity error;
    assert SOR = '1' report "Error in test case #1922/2803" severity error;
    assert SOL = '1' report "Error in test case #1922/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1923/2803" severity error;
    assert SOR = '1' report "Error in test case #1923/2803" severity error;
    assert SOL = '1' report "Error in test case #1923/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1924/2803" severity error;
    assert SOR = '1' report "Error in test case #1924/2803" severity error;
    assert SOL = '1' report "Error in test case #1924/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1925/2803" severity error;
    assert SOR = '1' report "Error in test case #1925/2803" severity error;
    assert SOL = '1' report "Error in test case #1925/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1926/2803" severity error;
    assert SOR = '1' report "Error in test case #1926/2803" severity error;
    assert SOL = '1' report "Error in test case #1926/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1927/2803" severity error;
    assert SOR = '1' report "Error in test case #1927/2803" severity error;
    assert SOL = '1' report "Error in test case #1927/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1928/2803" severity error;
    assert SOR = '1' report "Error in test case #1928/2803" severity error;
    assert SOL = '1' report "Error in test case #1928/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1929/2803" severity error;
    assert SOR = '1' report "Error in test case #1929/2803" severity error;
    assert SOL = '1' report "Error in test case #1929/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1930/2803" severity error;
    assert SOR = '1' report "Error in test case #1930/2803" severity error;
    assert SOL = '1' report "Error in test case #1930/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1931/2803" severity error;
    assert SOR = '1' report "Error in test case #1931/2803" severity error;
    assert SOL = '1' report "Error in test case #1931/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1932/2803" severity error;
    assert SOR = '1' report "Error in test case #1932/2803" severity error;
    assert SOL = '1' report "Error in test case #1932/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1933/2803" severity error;
    assert SOR = '1' report "Error in test case #1933/2803" severity error;
    assert SOL = '1' report "Error in test case #1933/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1934/2803" severity error;
    assert SOR = '1' report "Error in test case #1934/2803" severity error;
    assert SOL = '1' report "Error in test case #1934/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1935/2803" severity error;
    assert SOR = '1' report "Error in test case #1935/2803" severity error;
    assert SOL = '1' report "Error in test case #1935/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1936/2803" severity error;
    assert SOR = '1' report "Error in test case #1936/2803" severity error;
    assert SOL = '1' report "Error in test case #1936/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1937/2803" severity error;
    assert SOR = '1' report "Error in test case #1937/2803" severity error;
    assert SOL = '1' report "Error in test case #1937/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1938/2803" severity error;
    assert SOR = '1' report "Error in test case #1938/2803" severity error;
    assert SOL = '1' report "Error in test case #1938/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1939/2803" severity error;
    assert SOR = '1' report "Error in test case #1939/2803" severity error;
    assert SOL = '1' report "Error in test case #1939/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1940/2803" severity error;
    assert SOR = '1' report "Error in test case #1940/2803" severity error;
    assert SOL = '1' report "Error in test case #1940/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1941/2803" severity error;
    assert SOR = '1' report "Error in test case #1941/2803" severity error;
    assert SOL = '1' report "Error in test case #1941/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1942/2803" severity error;
    assert SOR = '1' report "Error in test case #1942/2803" severity error;
    assert SOL = '1' report "Error in test case #1942/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1943/2803" severity error;
    assert SOR = '1' report "Error in test case #1943/2803" severity error;
    assert SOL = '1' report "Error in test case #1943/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #1944/2803" severity error;
    assert SOR = '1' report "Error in test case #1944/2803" severity error;
    assert SOL = '1' report "Error in test case #1944/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1945/2803" severity error;
    assert SOR = '0' report "Error in test case #1945/2803" severity error;
    assert SOL = '0' report "Error in test case #1945/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1946/2803" severity error;
    assert SOR = '0' report "Error in test case #1946/2803" severity error;
    assert SOL = '0' report "Error in test case #1946/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1947/2803" severity error;
    assert SOR = '0' report "Error in test case #1947/2803" severity error;
    assert SOL = '0' report "Error in test case #1947/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1948/2803" severity error;
    assert SOR = '0' report "Error in test case #1948/2803" severity error;
    assert SOL = '0' report "Error in test case #1948/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1949/2803" severity error;
    assert SOR = '0' report "Error in test case #1949/2803" severity error;
    assert SOL = '0' report "Error in test case #1949/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1950/2803" severity error;
    assert SOR = '0' report "Error in test case #1950/2803" severity error;
    assert SOL = '0' report "Error in test case #1950/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1951/2803" severity error;
    assert SOR = '0' report "Error in test case #1951/2803" severity error;
    assert SOL = '0' report "Error in test case #1951/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1952/2803" severity error;
    assert SOR = '0' report "Error in test case #1952/2803" severity error;
    assert SOL = '0' report "Error in test case #1952/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1953/2803" severity error;
    assert SOR = '0' report "Error in test case #1953/2803" severity error;
    assert SOL = '0' report "Error in test case #1953/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1954/2803" severity error;
    assert SOR = '0' report "Error in test case #1954/2803" severity error;
    assert SOL = '0' report "Error in test case #1954/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1955/2803" severity error;
    assert SOR = '0' report "Error in test case #1955/2803" severity error;
    assert SOL = '0' report "Error in test case #1955/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1956/2803" severity error;
    assert SOR = '0' report "Error in test case #1956/2803" severity error;
    assert SOL = '0' report "Error in test case #1956/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1957/2803" severity error;
    assert SOR = '0' report "Error in test case #1957/2803" severity error;
    assert SOL = '0' report "Error in test case #1957/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1958/2803" severity error;
    assert SOR = '0' report "Error in test case #1958/2803" severity error;
    assert SOL = '0' report "Error in test case #1958/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1959/2803" severity error;
    assert SOR = '0' report "Error in test case #1959/2803" severity error;
    assert SOL = '0' report "Error in test case #1959/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1960/2803" severity error;
    assert SOR = '0' report "Error in test case #1960/2803" severity error;
    assert SOL = '0' report "Error in test case #1960/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1961/2803" severity error;
    assert SOR = '0' report "Error in test case #1961/2803" severity error;
    assert SOL = '0' report "Error in test case #1961/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1962/2803" severity error;
    assert SOR = '0' report "Error in test case #1962/2803" severity error;
    assert SOL = '0' report "Error in test case #1962/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1963/2803" severity error;
    assert SOR = '0' report "Error in test case #1963/2803" severity error;
    assert SOL = '0' report "Error in test case #1963/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1964/2803" severity error;
    assert SOR = '0' report "Error in test case #1964/2803" severity error;
    assert SOL = '0' report "Error in test case #1964/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1965/2803" severity error;
    assert SOR = '0' report "Error in test case #1965/2803" severity error;
    assert SOL = '0' report "Error in test case #1965/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1966/2803" severity error;
    assert SOR = '0' report "Error in test case #1966/2803" severity error;
    assert SOL = '0' report "Error in test case #1966/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1967/2803" severity error;
    assert SOR = '0' report "Error in test case #1967/2803" severity error;
    assert SOL = '0' report "Error in test case #1967/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1968/2803" severity error;
    assert SOR = '0' report "Error in test case #1968/2803" severity error;
    assert SOL = '0' report "Error in test case #1968/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1969/2803" severity error;
    assert SOR = '0' report "Error in test case #1969/2803" severity error;
    assert SOL = '0' report "Error in test case #1969/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1970/2803" severity error;
    assert SOR = '0' report "Error in test case #1970/2803" severity error;
    assert SOL = '0' report "Error in test case #1970/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1971/2803" severity error;
    assert SOR = '0' report "Error in test case #1971/2803" severity error;
    assert SOL = '0' report "Error in test case #1971/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1972/2803" severity error;
    assert SOR = '0' report "Error in test case #1972/2803" severity error;
    assert SOL = '0' report "Error in test case #1972/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1973/2803" severity error;
    assert SOR = '0' report "Error in test case #1973/2803" severity error;
    assert SOL = '0' report "Error in test case #1973/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1974/2803" severity error;
    assert SOR = '0' report "Error in test case #1974/2803" severity error;
    assert SOL = '0' report "Error in test case #1974/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1975/2803" severity error;
    assert SOR = '0' report "Error in test case #1975/2803" severity error;
    assert SOL = '0' report "Error in test case #1975/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1976/2803" severity error;
    assert SOR = '0' report "Error in test case #1976/2803" severity error;
    assert SOL = '0' report "Error in test case #1976/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1977/2803" severity error;
    assert SOR = '0' report "Error in test case #1977/2803" severity error;
    assert SOL = '0' report "Error in test case #1977/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1978/2803" severity error;
    assert SOR = '0' report "Error in test case #1978/2803" severity error;
    assert SOL = '0' report "Error in test case #1978/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1979/2803" severity error;
    assert SOR = '0' report "Error in test case #1979/2803" severity error;
    assert SOL = '0' report "Error in test case #1979/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1980/2803" severity error;
    assert SOR = '0' report "Error in test case #1980/2803" severity error;
    assert SOL = '0' report "Error in test case #1980/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1981/2803" severity error;
    assert SOR = '0' report "Error in test case #1981/2803" severity error;
    assert SOL = '0' report "Error in test case #1981/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1982/2803" severity error;
    assert SOR = '0' report "Error in test case #1982/2803" severity error;
    assert SOL = '0' report "Error in test case #1982/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1983/2803" severity error;
    assert SOR = '0' report "Error in test case #1983/2803" severity error;
    assert SOL = '0' report "Error in test case #1983/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1984/2803" severity error;
    assert SOR = '0' report "Error in test case #1984/2803" severity error;
    assert SOL = '0' report "Error in test case #1984/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1985/2803" severity error;
    assert SOR = '0' report "Error in test case #1985/2803" severity error;
    assert SOL = '0' report "Error in test case #1985/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1986/2803" severity error;
    assert SOR = '0' report "Error in test case #1986/2803" severity error;
    assert SOL = '0' report "Error in test case #1986/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1987/2803" severity error;
    assert SOR = '0' report "Error in test case #1987/2803" severity error;
    assert SOL = '0' report "Error in test case #1987/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1988/2803" severity error;
    assert SOR = '0' report "Error in test case #1988/2803" severity error;
    assert SOL = '0' report "Error in test case #1988/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1989/2803" severity error;
    assert SOR = '0' report "Error in test case #1989/2803" severity error;
    assert SOL = '0' report "Error in test case #1989/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1990/2803" severity error;
    assert SOR = '0' report "Error in test case #1990/2803" severity error;
    assert SOL = '0' report "Error in test case #1990/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1991/2803" severity error;
    assert SOR = '0' report "Error in test case #1991/2803" severity error;
    assert SOL = '0' report "Error in test case #1991/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1992/2803" severity error;
    assert SOR = '0' report "Error in test case #1992/2803" severity error;
    assert SOL = '0' report "Error in test case #1992/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1993/2803" severity error;
    assert SOR = '0' report "Error in test case #1993/2803" severity error;
    assert SOL = '0' report "Error in test case #1993/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1994/2803" severity error;
    assert SOR = '0' report "Error in test case #1994/2803" severity error;
    assert SOL = '0' report "Error in test case #1994/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1995/2803" severity error;
    assert SOR = '0' report "Error in test case #1995/2803" severity error;
    assert SOL = '0' report "Error in test case #1995/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1996/2803" severity error;
    assert SOR = '0' report "Error in test case #1996/2803" severity error;
    assert SOL = '0' report "Error in test case #1996/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1997/2803" severity error;
    assert SOR = '0' report "Error in test case #1997/2803" severity error;
    assert SOL = '0' report "Error in test case #1997/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1998/2803" severity error;
    assert SOR = '0' report "Error in test case #1998/2803" severity error;
    assert SOL = '0' report "Error in test case #1998/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #1999/2803" severity error;
    assert SOR = '0' report "Error in test case #1999/2803" severity error;
    assert SOL = '0' report "Error in test case #1999/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2000/2803" severity error;
    assert SOR = '0' report "Error in test case #2000/2803" severity error;
    assert SOL = '0' report "Error in test case #2000/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2001/2803" severity error;
    assert SOR = '0' report "Error in test case #2001/2803" severity error;
    assert SOL = '0' report "Error in test case #2001/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2002/2803" severity error;
    assert SOR = '0' report "Error in test case #2002/2803" severity error;
    assert SOL = '0' report "Error in test case #2002/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "100";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2003/2803" severity error;
    assert SOR = '0' report "Error in test case #2003/2803" severity error;
    assert SOL = '0' report "Error in test case #2003/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2004/2803" severity error;
    assert SOR = '0' report "Error in test case #2004/2803" severity error;
    assert SOL = '0' report "Error in test case #2004/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2005/2803" severity error;
    assert SOR = '0' report "Error in test case #2005/2803" severity error;
    assert SOL = '0' report "Error in test case #2005/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2006/2803" severity error;
    assert SOR = '0' report "Error in test case #2006/2803" severity error;
    assert SOL = '0' report "Error in test case #2006/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2007/2803" severity error;
    assert SOR = '0' report "Error in test case #2007/2803" severity error;
    assert SOL = '0' report "Error in test case #2007/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2008/2803" severity error;
    assert SOR = '0' report "Error in test case #2008/2803" severity error;
    assert SOL = '0' report "Error in test case #2008/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2009/2803" severity error;
    assert SOR = '0' report "Error in test case #2009/2803" severity error;
    assert SOL = '0' report "Error in test case #2009/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2010/2803" severity error;
    assert SOR = '0' report "Error in test case #2010/2803" severity error;
    assert SOL = '0' report "Error in test case #2010/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2011/2803" severity error;
    assert SOR = '0' report "Error in test case #2011/2803" severity error;
    assert SOL = '0' report "Error in test case #2011/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2012/2803" severity error;
    assert SOR = '0' report "Error in test case #2012/2803" severity error;
    assert SOL = '0' report "Error in test case #2012/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2013/2803" severity error;
    assert SOR = '0' report "Error in test case #2013/2803" severity error;
    assert SOL = '0' report "Error in test case #2013/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2014/2803" severity error;
    assert SOR = '0' report "Error in test case #2014/2803" severity error;
    assert SOL = '0' report "Error in test case #2014/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2015/2803" severity error;
    assert SOR = '0' report "Error in test case #2015/2803" severity error;
    assert SOL = '0' report "Error in test case #2015/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2016/2803" severity error;
    assert SOR = '0' report "Error in test case #2016/2803" severity error;
    assert SOL = '0' report "Error in test case #2016/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2017/2803" severity error;
    assert SOR = '0' report "Error in test case #2017/2803" severity error;
    assert SOL = '0' report "Error in test case #2017/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2018/2803" severity error;
    assert SOR = '0' report "Error in test case #2018/2803" severity error;
    assert SOL = '0' report "Error in test case #2018/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2019/2803" severity error;
    assert SOR = '0' report "Error in test case #2019/2803" severity error;
    assert SOL = '0' report "Error in test case #2019/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2020/2803" severity error;
    assert SOR = '0' report "Error in test case #2020/2803" severity error;
    assert SOL = '0' report "Error in test case #2020/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2021/2803" severity error;
    assert SOR = '0' report "Error in test case #2021/2803" severity error;
    assert SOL = '0' report "Error in test case #2021/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2022/2803" severity error;
    assert SOR = '0' report "Error in test case #2022/2803" severity error;
    assert SOL = '0' report "Error in test case #2022/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2023/2803" severity error;
    assert SOR = '0' report "Error in test case #2023/2803" severity error;
    assert SOL = '0' report "Error in test case #2023/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2024/2803" severity error;
    assert SOR = '0' report "Error in test case #2024/2803" severity error;
    assert SOL = '0' report "Error in test case #2024/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2025/2803" severity error;
    assert SOR = '0' report "Error in test case #2025/2803" severity error;
    assert SOL = '0' report "Error in test case #2025/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2026/2803" severity error;
    assert SOR = '0' report "Error in test case #2026/2803" severity error;
    assert SOL = '0' report "Error in test case #2026/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2027/2803" severity error;
    assert SOR = '0' report "Error in test case #2027/2803" severity error;
    assert SOL = '0' report "Error in test case #2027/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2028/2803" severity error;
    assert SOR = '0' report "Error in test case #2028/2803" severity error;
    assert SOL = '0' report "Error in test case #2028/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2029/2803" severity error;
    assert SOR = '0' report "Error in test case #2029/2803" severity error;
    assert SOL = '0' report "Error in test case #2029/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2030/2803" severity error;
    assert SOR = '0' report "Error in test case #2030/2803" severity error;
    assert SOL = '0' report "Error in test case #2030/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2031/2803" severity error;
    assert SOR = '0' report "Error in test case #2031/2803" severity error;
    assert SOL = '0' report "Error in test case #2031/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2032/2803" severity error;
    assert SOR = '0' report "Error in test case #2032/2803" severity error;
    assert SOL = '0' report "Error in test case #2032/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2033/2803" severity error;
    assert SOR = '0' report "Error in test case #2033/2803" severity error;
    assert SOL = '0' report "Error in test case #2033/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2034/2803" severity error;
    assert SOR = '0' report "Error in test case #2034/2803" severity error;
    assert SOL = '0' report "Error in test case #2034/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2035/2803" severity error;
    assert SOR = '0' report "Error in test case #2035/2803" severity error;
    assert SOL = '0' report "Error in test case #2035/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2036/2803" severity error;
    assert SOR = '0' report "Error in test case #2036/2803" severity error;
    assert SOL = '0' report "Error in test case #2036/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2037/2803" severity error;
    assert SOR = '0' report "Error in test case #2037/2803" severity error;
    assert SOL = '0' report "Error in test case #2037/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2038/2803" severity error;
    assert SOR = '0' report "Error in test case #2038/2803" severity error;
    assert SOL = '0' report "Error in test case #2038/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2039/2803" severity error;
    assert SOR = '0' report "Error in test case #2039/2803" severity error;
    assert SOL = '0' report "Error in test case #2039/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2040/2803" severity error;
    assert SOR = '0' report "Error in test case #2040/2803" severity error;
    assert SOL = '0' report "Error in test case #2040/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2041/2803" severity error;
    assert SOR = '0' report "Error in test case #2041/2803" severity error;
    assert SOL = '0' report "Error in test case #2041/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2042/2803" severity error;
    assert SOR = '0' report "Error in test case #2042/2803" severity error;
    assert SOL = '0' report "Error in test case #2042/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2043/2803" severity error;
    assert SOR = '0' report "Error in test case #2043/2803" severity error;
    assert SOL = '0' report "Error in test case #2043/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2044/2803" severity error;
    assert SOR = '0' report "Error in test case #2044/2803" severity error;
    assert SOL = '0' report "Error in test case #2044/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2045/2803" severity error;
    assert SOR = '0' report "Error in test case #2045/2803" severity error;
    assert SOL = '0' report "Error in test case #2045/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2046/2803" severity error;
    assert SOR = '0' report "Error in test case #2046/2803" severity error;
    assert SOL = '0' report "Error in test case #2046/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2047/2803" severity error;
    assert SOR = '0' report "Error in test case #2047/2803" severity error;
    assert SOL = '0' report "Error in test case #2047/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2048/2803" severity error;
    assert SOR = '0' report "Error in test case #2048/2803" severity error;
    assert SOL = '0' report "Error in test case #2048/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2049/2803" severity error;
    assert SOR = '0' report "Error in test case #2049/2803" severity error;
    assert SOL = '0' report "Error in test case #2049/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2050/2803" severity error;
    assert SOR = '0' report "Error in test case #2050/2803" severity error;
    assert SOL = '0' report "Error in test case #2050/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2051/2803" severity error;
    assert SOR = '0' report "Error in test case #2051/2803" severity error;
    assert SOL = '0' report "Error in test case #2051/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2052/2803" severity error;
    assert SOR = '0' report "Error in test case #2052/2803" severity error;
    assert SOL = '0' report "Error in test case #2052/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2053/2803" severity error;
    assert SOR = '0' report "Error in test case #2053/2803" severity error;
    assert SOL = '0' report "Error in test case #2053/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2054/2803" severity error;
    assert SOR = '0' report "Error in test case #2054/2803" severity error;
    assert SOL = '0' report "Error in test case #2054/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2055/2803" severity error;
    assert SOR = '0' report "Error in test case #2055/2803" severity error;
    assert SOL = '0' report "Error in test case #2055/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2056/2803" severity error;
    assert SOR = '0' report "Error in test case #2056/2803" severity error;
    assert SOL = '0' report "Error in test case #2056/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2057/2803" severity error;
    assert SOR = '0' report "Error in test case #2057/2803" severity error;
    assert SOL = '0' report "Error in test case #2057/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2058/2803" severity error;
    assert SOR = '0' report "Error in test case #2058/2803" severity error;
    assert SOL = '0' report "Error in test case #2058/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2059/2803" severity error;
    assert SOR = '0' report "Error in test case #2059/2803" severity error;
    assert SOL = '0' report "Error in test case #2059/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2060/2803" severity error;
    assert SOR = '0' report "Error in test case #2060/2803" severity error;
    assert SOL = '0' report "Error in test case #2060/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2061/2803" severity error;
    assert SOR = '0' report "Error in test case #2061/2803" severity error;
    assert SOL = '0' report "Error in test case #2061/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2062/2803" severity error;
    assert SOR = '0' report "Error in test case #2062/2803" severity error;
    assert SOL = '0' report "Error in test case #2062/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2063/2803" severity error;
    assert SOR = '0' report "Error in test case #2063/2803" severity error;
    assert SOL = '0' report "Error in test case #2063/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2064/2803" severity error;
    assert SOR = '0' report "Error in test case #2064/2803" severity error;
    assert SOL = '0' report "Error in test case #2064/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2065/2803" severity error;
    assert SOR = '0' report "Error in test case #2065/2803" severity error;
    assert SOL = '0' report "Error in test case #2065/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2066/2803" severity error;
    assert SOR = '0' report "Error in test case #2066/2803" severity error;
    assert SOL = '0' report "Error in test case #2066/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2067/2803" severity error;
    assert SOR = '0' report "Error in test case #2067/2803" severity error;
    assert SOL = '0' report "Error in test case #2067/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2068/2803" severity error;
    assert SOR = '0' report "Error in test case #2068/2803" severity error;
    assert SOL = '0' report "Error in test case #2068/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2069/2803" severity error;
    assert SOR = '0' report "Error in test case #2069/2803" severity error;
    assert SOL = '0' report "Error in test case #2069/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2070/2803" severity error;
    assert SOR = '0' report "Error in test case #2070/2803" severity error;
    assert SOL = '0' report "Error in test case #2070/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2071/2803" severity error;
    assert SOR = '0' report "Error in test case #2071/2803" severity error;
    assert SOL = '0' report "Error in test case #2071/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2072/2803" severity error;
    assert SOR = '0' report "Error in test case #2072/2803" severity error;
    assert SOL = '0' report "Error in test case #2072/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2073/2803" severity error;
    assert SOR = '0' report "Error in test case #2073/2803" severity error;
    assert SOL = '0' report "Error in test case #2073/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2074/2803" severity error;
    assert SOR = '0' report "Error in test case #2074/2803" severity error;
    assert SOL = '0' report "Error in test case #2074/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2075/2803" severity error;
    assert SOR = '0' report "Error in test case #2075/2803" severity error;
    assert SOL = '0' report "Error in test case #2075/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2076/2803" severity error;
    assert SOR = '0' report "Error in test case #2076/2803" severity error;
    assert SOL = '0' report "Error in test case #2076/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2077/2803" severity error;
    assert SOR = '0' report "Error in test case #2077/2803" severity error;
    assert SOL = '0' report "Error in test case #2077/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2078/2803" severity error;
    assert SOR = '0' report "Error in test case #2078/2803" severity error;
    assert SOL = '0' report "Error in test case #2078/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2079/2803" severity error;
    assert SOR = '0' report "Error in test case #2079/2803" severity error;
    assert SOL = '0' report "Error in test case #2079/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2080/2803" severity error;
    assert SOR = '0' report "Error in test case #2080/2803" severity error;
    assert SOL = '0' report "Error in test case #2080/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2081/2803" severity error;
    assert SOR = '0' report "Error in test case #2081/2803" severity error;
    assert SOL = '0' report "Error in test case #2081/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2082/2803" severity error;
    assert SOR = '0' report "Error in test case #2082/2803" severity error;
    assert SOL = '0' report "Error in test case #2082/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2083/2803" severity error;
    assert SOR = '0' report "Error in test case #2083/2803" severity error;
    assert SOL = '0' report "Error in test case #2083/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2084/2803" severity error;
    assert SOR = '0' report "Error in test case #2084/2803" severity error;
    assert SOL = '0' report "Error in test case #2084/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2085/2803" severity error;
    assert SOR = '0' report "Error in test case #2085/2803" severity error;
    assert SOL = '0' report "Error in test case #2085/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2086/2803" severity error;
    assert SOR = '0' report "Error in test case #2086/2803" severity error;
    assert SOL = '0' report "Error in test case #2086/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2087/2803" severity error;
    assert SOR = '0' report "Error in test case #2087/2803" severity error;
    assert SOL = '0' report "Error in test case #2087/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2088/2803" severity error;
    assert SOR = '0' report "Error in test case #2088/2803" severity error;
    assert SOL = '0' report "Error in test case #2088/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2089/2803" severity error;
    assert SOR = '0' report "Error in test case #2089/2803" severity error;
    assert SOL = '0' report "Error in test case #2089/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2090/2803" severity error;
    assert SOR = '0' report "Error in test case #2090/2803" severity error;
    assert SOL = '0' report "Error in test case #2090/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2091/2803" severity error;
    assert SOR = '0' report "Error in test case #2091/2803" severity error;
    assert SOL = '0' report "Error in test case #2091/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2092/2803" severity error;
    assert SOR = '0' report "Error in test case #2092/2803" severity error;
    assert SOL = '0' report "Error in test case #2092/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2093/2803" severity error;
    assert SOR = '0' report "Error in test case #2093/2803" severity error;
    assert SOL = '0' report "Error in test case #2093/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2094/2803" severity error;
    assert SOR = '0' report "Error in test case #2094/2803" severity error;
    assert SOL = '0' report "Error in test case #2094/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2095/2803" severity error;
    assert SOR = '0' report "Error in test case #2095/2803" severity error;
    assert SOL = '0' report "Error in test case #2095/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2096/2803" severity error;
    assert SOR = '0' report "Error in test case #2096/2803" severity error;
    assert SOL = '0' report "Error in test case #2096/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2097/2803" severity error;
    assert SOR = '0' report "Error in test case #2097/2803" severity error;
    assert SOL = '0' report "Error in test case #2097/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2098/2803" severity error;
    assert SOR = '0' report "Error in test case #2098/2803" severity error;
    assert SOL = '0' report "Error in test case #2098/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2099/2803" severity error;
    assert SOR = '0' report "Error in test case #2099/2803" severity error;
    assert SOL = '0' report "Error in test case #2099/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2100/2803" severity error;
    assert SOR = '0' report "Error in test case #2100/2803" severity error;
    assert SOL = '0' report "Error in test case #2100/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2101/2803" severity error;
    assert SOR = '0' report "Error in test case #2101/2803" severity error;
    assert SOL = '0' report "Error in test case #2101/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2102/2803" severity error;
    assert SOR = '0' report "Error in test case #2102/2803" severity error;
    assert SOL = '0' report "Error in test case #2102/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2103/2803" severity error;
    assert SOR = '0' report "Error in test case #2103/2803" severity error;
    assert SOL = '0' report "Error in test case #2103/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2104/2803" severity error;
    assert SOR = '0' report "Error in test case #2104/2803" severity error;
    assert SOL = '0' report "Error in test case #2104/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2105/2803" severity error;
    assert SOR = '0' report "Error in test case #2105/2803" severity error;
    assert SOL = '0' report "Error in test case #2105/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2106/2803" severity error;
    assert SOR = '0' report "Error in test case #2106/2803" severity error;
    assert SOL = '0' report "Error in test case #2106/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2107/2803" severity error;
    assert SOR = '0' report "Error in test case #2107/2803" severity error;
    assert SOL = '0' report "Error in test case #2107/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2108/2803" severity error;
    assert SOR = '0' report "Error in test case #2108/2803" severity error;
    assert SOL = '0' report "Error in test case #2108/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2109/2803" severity error;
    assert SOR = '0' report "Error in test case #2109/2803" severity error;
    assert SOL = '0' report "Error in test case #2109/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2110/2803" severity error;
    assert SOR = '0' report "Error in test case #2110/2803" severity error;
    assert SOL = '0' report "Error in test case #2110/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2111/2803" severity error;
    assert SOR = '0' report "Error in test case #2111/2803" severity error;
    assert SOL = '0' report "Error in test case #2111/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2112/2803" severity error;
    assert SOR = '0' report "Error in test case #2112/2803" severity error;
    assert SOL = '0' report "Error in test case #2112/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2113/2803" severity error;
    assert SOR = '0' report "Error in test case #2113/2803" severity error;
    assert SOL = '0' report "Error in test case #2113/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2114/2803" severity error;
    assert SOR = '0' report "Error in test case #2114/2803" severity error;
    assert SOL = '0' report "Error in test case #2114/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2115/2803" severity error;
    assert SOR = '0' report "Error in test case #2115/2803" severity error;
    assert SOL = '0' report "Error in test case #2115/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2116/2803" severity error;
    assert SOR = '0' report "Error in test case #2116/2803" severity error;
    assert SOL = '0' report "Error in test case #2116/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2117/2803" severity error;
    assert SOR = '0' report "Error in test case #2117/2803" severity error;
    assert SOL = '0' report "Error in test case #2117/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2118/2803" severity error;
    assert SOR = '0' report "Error in test case #2118/2803" severity error;
    assert SOL = '0' report "Error in test case #2118/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2119/2803" severity error;
    assert SOR = '0' report "Error in test case #2119/2803" severity error;
    assert SOL = '0' report "Error in test case #2119/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2120/2803" severity error;
    assert SOR = '0' report "Error in test case #2120/2803" severity error;
    assert SOL = '0' report "Error in test case #2120/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2121/2803" severity error;
    assert SOR = '0' report "Error in test case #2121/2803" severity error;
    assert SOL = '0' report "Error in test case #2121/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2122/2803" severity error;
    assert SOR = '0' report "Error in test case #2122/2803" severity error;
    assert SOL = '0' report "Error in test case #2122/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2123/2803" severity error;
    assert SOR = '0' report "Error in test case #2123/2803" severity error;
    assert SOL = '0' report "Error in test case #2123/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2124/2803" severity error;
    assert SOR = '0' report "Error in test case #2124/2803" severity error;
    assert SOL = '0' report "Error in test case #2124/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2125/2803" severity error;
    assert SOR = '0' report "Error in test case #2125/2803" severity error;
    assert SOL = '0' report "Error in test case #2125/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2126/2803" severity error;
    assert SOR = '0' report "Error in test case #2126/2803" severity error;
    assert SOL = '0' report "Error in test case #2126/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2127/2803" severity error;
    assert SOR = '0' report "Error in test case #2127/2803" severity error;
    assert SOL = '0' report "Error in test case #2127/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2128/2803" severity error;
    assert SOR = '0' report "Error in test case #2128/2803" severity error;
    assert SOL = '0' report "Error in test case #2128/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2129/2803" severity error;
    assert SOR = '0' report "Error in test case #2129/2803" severity error;
    assert SOL = '0' report "Error in test case #2129/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2130/2803" severity error;
    assert SOR = '0' report "Error in test case #2130/2803" severity error;
    assert SOL = '0' report "Error in test case #2130/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2131/2803" severity error;
    assert SOR = '0' report "Error in test case #2131/2803" severity error;
    assert SOL = '0' report "Error in test case #2131/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2132/2803" severity error;
    assert SOR = '0' report "Error in test case #2132/2803" severity error;
    assert SOL = '0' report "Error in test case #2132/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2133/2803" severity error;
    assert SOR = '0' report "Error in test case #2133/2803" severity error;
    assert SOL = '0' report "Error in test case #2133/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2134/2803" severity error;
    assert SOR = '0' report "Error in test case #2134/2803" severity error;
    assert SOL = '0' report "Error in test case #2134/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2135/2803" severity error;
    assert SOR = '0' report "Error in test case #2135/2803" severity error;
    assert SOL = '0' report "Error in test case #2135/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2136/2803" severity error;
    assert SOR = '0' report "Error in test case #2136/2803" severity error;
    assert SOL = '0' report "Error in test case #2136/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2137/2803" severity error;
    assert SOR = '0' report "Error in test case #2137/2803" severity error;
    assert SOL = '0' report "Error in test case #2137/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2138/2803" severity error;
    assert SOR = '0' report "Error in test case #2138/2803" severity error;
    assert SOL = '0' report "Error in test case #2138/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2139/2803" severity error;
    assert SOR = '0' report "Error in test case #2139/2803" severity error;
    assert SOL = '0' report "Error in test case #2139/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2140/2803" severity error;
    assert SOR = '0' report "Error in test case #2140/2803" severity error;
    assert SOL = '0' report "Error in test case #2140/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2141/2803" severity error;
    assert SOR = '0' report "Error in test case #2141/2803" severity error;
    assert SOL = '0' report "Error in test case #2141/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2142/2803" severity error;
    assert SOR = '0' report "Error in test case #2142/2803" severity error;
    assert SOL = '0' report "Error in test case #2142/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2143/2803" severity error;
    assert SOR = '0' report "Error in test case #2143/2803" severity error;
    assert SOL = '0' report "Error in test case #2143/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2144/2803" severity error;
    assert SOR = '0' report "Error in test case #2144/2803" severity error;
    assert SOL = '0' report "Error in test case #2144/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2145/2803" severity error;
    assert SOR = '0' report "Error in test case #2145/2803" severity error;
    assert SOL = '0' report "Error in test case #2145/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2146/2803" severity error;
    assert SOR = '0' report "Error in test case #2146/2803" severity error;
    assert SOL = '0' report "Error in test case #2146/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2147/2803" severity error;
    assert SOR = '0' report "Error in test case #2147/2803" severity error;
    assert SOL = '0' report "Error in test case #2147/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2148/2803" severity error;
    assert SOR = '0' report "Error in test case #2148/2803" severity error;
    assert SOL = '0' report "Error in test case #2148/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2149/2803" severity error;
    assert SOR = '0' report "Error in test case #2149/2803" severity error;
    assert SOL = '0' report "Error in test case #2149/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2150/2803" severity error;
    assert SOR = '0' report "Error in test case #2150/2803" severity error;
    assert SOL = '0' report "Error in test case #2150/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2151/2803" severity error;
    assert SOR = '0' report "Error in test case #2151/2803" severity error;
    assert SOL = '0' report "Error in test case #2151/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2152/2803" severity error;
    assert SOR = '0' report "Error in test case #2152/2803" severity error;
    assert SOL = '0' report "Error in test case #2152/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2153/2803" severity error;
    assert SOR = '0' report "Error in test case #2153/2803" severity error;
    assert SOL = '0' report "Error in test case #2153/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2154/2803" severity error;
    assert SOR = '0' report "Error in test case #2154/2803" severity error;
    assert SOL = '0' report "Error in test case #2154/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2155/2803" severity error;
    assert SOR = '0' report "Error in test case #2155/2803" severity error;
    assert SOL = '0' report "Error in test case #2155/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2156/2803" severity error;
    assert SOR = '0' report "Error in test case #2156/2803" severity error;
    assert SOL = '0' report "Error in test case #2156/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2157/2803" severity error;
    assert SOR = '0' report "Error in test case #2157/2803" severity error;
    assert SOL = '0' report "Error in test case #2157/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2158/2803" severity error;
    assert SOR = '0' report "Error in test case #2158/2803" severity error;
    assert SOL = '0' report "Error in test case #2158/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2159/2803" severity error;
    assert SOR = '0' report "Error in test case #2159/2803" severity error;
    assert SOL = '0' report "Error in test case #2159/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2160/2803" severity error;
    assert SOR = '0' report "Error in test case #2160/2803" severity error;
    assert SOL = '0' report "Error in test case #2160/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2161/2803" severity error;
    assert SOR = '0' report "Error in test case #2161/2803" severity error;
    assert SOL = '0' report "Error in test case #2161/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2162/2803" severity error;
    assert SOR = '0' report "Error in test case #2162/2803" severity error;
    assert SOL = '0' report "Error in test case #2162/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2163/2803" severity error;
    assert SOR = '0' report "Error in test case #2163/2803" severity error;
    assert SOL = '0' report "Error in test case #2163/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2164/2803" severity error;
    assert SOR = '0' report "Error in test case #2164/2803" severity error;
    assert SOL = '0' report "Error in test case #2164/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2165/2803" severity error;
    assert SOR = '0' report "Error in test case #2165/2803" severity error;
    assert SOL = '0' report "Error in test case #2165/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2166/2803" severity error;
    assert SOR = '0' report "Error in test case #2166/2803" severity error;
    assert SOL = '0' report "Error in test case #2166/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2167/2803" severity error;
    assert SOR = '0' report "Error in test case #2167/2803" severity error;
    assert SOL = '0' report "Error in test case #2167/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2168/2803" severity error;
    assert SOR = '0' report "Error in test case #2168/2803" severity error;
    assert SOL = '0' report "Error in test case #2168/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2169/2803" severity error;
    assert SOR = '0' report "Error in test case #2169/2803" severity error;
    assert SOL = '0' report "Error in test case #2169/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2170/2803" severity error;
    assert SOR = '0' report "Error in test case #2170/2803" severity error;
    assert SOL = '0' report "Error in test case #2170/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2171/2803" severity error;
    assert SOR = '0' report "Error in test case #2171/2803" severity error;
    assert SOL = '0' report "Error in test case #2171/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2172/2803" severity error;
    assert SOR = '0' report "Error in test case #2172/2803" severity error;
    assert SOL = '0' report "Error in test case #2172/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2173/2803" severity error;
    assert SOR = '0' report "Error in test case #2173/2803" severity error;
    assert SOL = '0' report "Error in test case #2173/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2174/2803" severity error;
    assert SOR = '0' report "Error in test case #2174/2803" severity error;
    assert SOL = '0' report "Error in test case #2174/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2175/2803" severity error;
    assert SOR = '0' report "Error in test case #2175/2803" severity error;
    assert SOL = '0' report "Error in test case #2175/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2176/2803" severity error;
    assert SOR = '0' report "Error in test case #2176/2803" severity error;
    assert SOL = '0' report "Error in test case #2176/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2177/2803" severity error;
    assert SOR = '0' report "Error in test case #2177/2803" severity error;
    assert SOL = '0' report "Error in test case #2177/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2178/2803" severity error;
    assert SOR = '0' report "Error in test case #2178/2803" severity error;
    assert SOL = '0' report "Error in test case #2178/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2179/2803" severity error;
    assert SOR = '0' report "Error in test case #2179/2803" severity error;
    assert SOL = '0' report "Error in test case #2179/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2180/2803" severity error;
    assert SOR = '0' report "Error in test case #2180/2803" severity error;
    assert SOL = '0' report "Error in test case #2180/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2181/2803" severity error;
    assert SOR = '0' report "Error in test case #2181/2803" severity error;
    assert SOL = '0' report "Error in test case #2181/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2182/2803" severity error;
    assert SOR = '0' report "Error in test case #2182/2803" severity error;
    assert SOL = '0' report "Error in test case #2182/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2183/2803" severity error;
    assert SOR = '0' report "Error in test case #2183/2803" severity error;
    assert SOL = '0' report "Error in test case #2183/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2184/2803" severity error;
    assert SOR = '0' report "Error in test case #2184/2803" severity error;
    assert SOL = '0' report "Error in test case #2184/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2185/2803" severity error;
    assert SOR = '0' report "Error in test case #2185/2803" severity error;
    assert SOL = '0' report "Error in test case #2185/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2186/2803" severity error;
    assert SOR = '0' report "Error in test case #2186/2803" severity error;
    assert SOL = '0' report "Error in test case #2186/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2187/2803" severity error;
    assert SOR = '0' report "Error in test case #2187/2803" severity error;
    assert SOL = '0' report "Error in test case #2187/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2188/2803" severity error;
    assert SOR = '0' report "Error in test case #2188/2803" severity error;
    assert SOL = '0' report "Error in test case #2188/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2189/2803" severity error;
    assert SOR = '0' report "Error in test case #2189/2803" severity error;
    assert SOL = '0' report "Error in test case #2189/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2190/2803" severity error;
    assert SOR = '0' report "Error in test case #2190/2803" severity error;
    assert SOL = '0' report "Error in test case #2190/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2191/2803" severity error;
    assert SOR = '0' report "Error in test case #2191/2803" severity error;
    assert SOL = '0' report "Error in test case #2191/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2192/2803" severity error;
    assert SOR = '0' report "Error in test case #2192/2803" severity error;
    assert SOL = '0' report "Error in test case #2192/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2193/2803" severity error;
    assert SOR = '0' report "Error in test case #2193/2803" severity error;
    assert SOL = '0' report "Error in test case #2193/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2194/2803" severity error;
    assert SOR = '0' report "Error in test case #2194/2803" severity error;
    assert SOL = '0' report "Error in test case #2194/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2195/2803" severity error;
    assert SOR = '0' report "Error in test case #2195/2803" severity error;
    assert SOL = '0' report "Error in test case #2195/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2196/2803" severity error;
    assert SOR = '0' report "Error in test case #2196/2803" severity error;
    assert SOL = '0' report "Error in test case #2196/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2197/2803" severity error;
    assert SOR = '0' report "Error in test case #2197/2803" severity error;
    assert SOL = '0' report "Error in test case #2197/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2198/2803" severity error;
    assert SOR = '0' report "Error in test case #2198/2803" severity error;
    assert SOL = '0' report "Error in test case #2198/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2199/2803" severity error;
    assert SOR = '0' report "Error in test case #2199/2803" severity error;
    assert SOL = '0' report "Error in test case #2199/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2200/2803" severity error;
    assert SOR = '0' report "Error in test case #2200/2803" severity error;
    assert SOL = '0' report "Error in test case #2200/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2201/2803" severity error;
    assert SOR = '0' report "Error in test case #2201/2803" severity error;
    assert SOL = '0' report "Error in test case #2201/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2202/2803" severity error;
    assert SOR = '0' report "Error in test case #2202/2803" severity error;
    assert SOL = '0' report "Error in test case #2202/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2203/2803" severity error;
    assert SOR = '0' report "Error in test case #2203/2803" severity error;
    assert SOL = '0' report "Error in test case #2203/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2204/2803" severity error;
    assert SOR = '0' report "Error in test case #2204/2803" severity error;
    assert SOL = '0' report "Error in test case #2204/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2205/2803" severity error;
    assert SOR = '0' report "Error in test case #2205/2803" severity error;
    assert SOL = '0' report "Error in test case #2205/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2206/2803" severity error;
    assert SOR = '0' report "Error in test case #2206/2803" severity error;
    assert SOL = '0' report "Error in test case #2206/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2207/2803" severity error;
    assert SOR = '0' report "Error in test case #2207/2803" severity error;
    assert SOL = '0' report "Error in test case #2207/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2208/2803" severity error;
    assert SOR = '0' report "Error in test case #2208/2803" severity error;
    assert SOL = '0' report "Error in test case #2208/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2209/2803" severity error;
    assert SOR = '0' report "Error in test case #2209/2803" severity error;
    assert SOL = '0' report "Error in test case #2209/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2210/2803" severity error;
    assert SOR = '0' report "Error in test case #2210/2803" severity error;
    assert SOL = '0' report "Error in test case #2210/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2211/2803" severity error;
    assert SOR = '0' report "Error in test case #2211/2803" severity error;
    assert SOL = '0' report "Error in test case #2211/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2212/2803" severity error;
    assert SOR = '0' report "Error in test case #2212/2803" severity error;
    assert SOL = '0' report "Error in test case #2212/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2213/2803" severity error;
    assert SOR = '0' report "Error in test case #2213/2803" severity error;
    assert SOL = '0' report "Error in test case #2213/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2214/2803" severity error;
    assert SOR = '0' report "Error in test case #2214/2803" severity error;
    assert SOL = '0' report "Error in test case #2214/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2215/2803" severity error;
    assert SOR = '0' report "Error in test case #2215/2803" severity error;
    assert SOL = '0' report "Error in test case #2215/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2216/2803" severity error;
    assert SOR = '0' report "Error in test case #2216/2803" severity error;
    assert SOL = '0' report "Error in test case #2216/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2217/2803" severity error;
    assert SOR = '0' report "Error in test case #2217/2803" severity error;
    assert SOL = '0' report "Error in test case #2217/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2218/2803" severity error;
    assert SOR = '0' report "Error in test case #2218/2803" severity error;
    assert SOL = '0' report "Error in test case #2218/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2219/2803" severity error;
    assert SOR = '0' report "Error in test case #2219/2803" severity error;
    assert SOL = '0' report "Error in test case #2219/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2220/2803" severity error;
    assert SOR = '0' report "Error in test case #2220/2803" severity error;
    assert SOL = '0' report "Error in test case #2220/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2221/2803" severity error;
    assert SOR = '0' report "Error in test case #2221/2803" severity error;
    assert SOL = '0' report "Error in test case #2221/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2222/2803" severity error;
    assert SOR = '0' report "Error in test case #2222/2803" severity error;
    assert SOL = '0' report "Error in test case #2222/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2223/2803" severity error;
    assert SOR = '0' report "Error in test case #2223/2803" severity error;
    assert SOL = '0' report "Error in test case #2223/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2224/2803" severity error;
    assert SOR = '0' report "Error in test case #2224/2803" severity error;
    assert SOL = '0' report "Error in test case #2224/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2225/2803" severity error;
    assert SOR = '0' report "Error in test case #2225/2803" severity error;
    assert SOL = '0' report "Error in test case #2225/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2226/2803" severity error;
    assert SOR = '0' report "Error in test case #2226/2803" severity error;
    assert SOL = '0' report "Error in test case #2226/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2227/2803" severity error;
    assert SOR = '0' report "Error in test case #2227/2803" severity error;
    assert SOL = '0' report "Error in test case #2227/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2228/2803" severity error;
    assert SOR = '0' report "Error in test case #2228/2803" severity error;
    assert SOL = '0' report "Error in test case #2228/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2229/2803" severity error;
    assert SOR = '0' report "Error in test case #2229/2803" severity error;
    assert SOL = '0' report "Error in test case #2229/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2230/2803" severity error;
    assert SOR = '0' report "Error in test case #2230/2803" severity error;
    assert SOL = '0' report "Error in test case #2230/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2231/2803" severity error;
    assert SOR = '0' report "Error in test case #2231/2803" severity error;
    assert SOL = '0' report "Error in test case #2231/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2232/2803" severity error;
    assert SOR = '0' report "Error in test case #2232/2803" severity error;
    assert SOL = '0' report "Error in test case #2232/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2233/2803" severity error;
    assert SOR = '0' report "Error in test case #2233/2803" severity error;
    assert SOL = '0' report "Error in test case #2233/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2234/2803" severity error;
    assert SOR = '0' report "Error in test case #2234/2803" severity error;
    assert SOL = '0' report "Error in test case #2234/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2235/2803" severity error;
    assert SOR = '0' report "Error in test case #2235/2803" severity error;
    assert SOL = '0' report "Error in test case #2235/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2236/2803" severity error;
    assert SOR = '0' report "Error in test case #2236/2803" severity error;
    assert SOL = '0' report "Error in test case #2236/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2237/2803" severity error;
    assert SOR = '0' report "Error in test case #2237/2803" severity error;
    assert SOL = '0' report "Error in test case #2237/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2238/2803" severity error;
    assert SOR = '0' report "Error in test case #2238/2803" severity error;
    assert SOL = '0' report "Error in test case #2238/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2239/2803" severity error;
    assert SOR = '0' report "Error in test case #2239/2803" severity error;
    assert SOL = '0' report "Error in test case #2239/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2240/2803" severity error;
    assert SOR = '0' report "Error in test case #2240/2803" severity error;
    assert SOL = '0' report "Error in test case #2240/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2241/2803" severity error;
    assert SOR = '0' report "Error in test case #2241/2803" severity error;
    assert SOL = '0' report "Error in test case #2241/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2242/2803" severity error;
    assert SOR = '0' report "Error in test case #2242/2803" severity error;
    assert SOL = '0' report "Error in test case #2242/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2243/2803" severity error;
    assert SOR = '0' report "Error in test case #2243/2803" severity error;
    assert SOL = '0' report "Error in test case #2243/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2244/2803" severity error;
    assert SOR = '0' report "Error in test case #2244/2803" severity error;
    assert SOL = '0' report "Error in test case #2244/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2245/2803" severity error;
    assert SOR = '0' report "Error in test case #2245/2803" severity error;
    assert SOL = '0' report "Error in test case #2245/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2246/2803" severity error;
    assert SOR = '0' report "Error in test case #2246/2803" severity error;
    assert SOL = '0' report "Error in test case #2246/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2247/2803" severity error;
    assert SOR = '0' report "Error in test case #2247/2803" severity error;
    assert SOL = '0' report "Error in test case #2247/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2248/2803" severity error;
    assert SOR = '0' report "Error in test case #2248/2803" severity error;
    assert SOL = '0' report "Error in test case #2248/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2249/2803" severity error;
    assert SOR = '0' report "Error in test case #2249/2803" severity error;
    assert SOL = '0' report "Error in test case #2249/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2250/2803" severity error;
    assert SOR = '0' report "Error in test case #2250/2803" severity error;
    assert SOL = '0' report "Error in test case #2250/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2251/2803" severity error;
    assert SOR = '0' report "Error in test case #2251/2803" severity error;
    assert SOL = '0' report "Error in test case #2251/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2252/2803" severity error;
    assert SOR = '0' report "Error in test case #2252/2803" severity error;
    assert SOL = '0' report "Error in test case #2252/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2253/2803" severity error;
    assert SOR = '0' report "Error in test case #2253/2803" severity error;
    assert SOL = '0' report "Error in test case #2253/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2254/2803" severity error;
    assert SOR = '0' report "Error in test case #2254/2803" severity error;
    assert SOL = '0' report "Error in test case #2254/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2255/2803" severity error;
    assert SOR = '0' report "Error in test case #2255/2803" severity error;
    assert SOL = '0' report "Error in test case #2255/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2256/2803" severity error;
    assert SOR = '0' report "Error in test case #2256/2803" severity error;
    assert SOL = '0' report "Error in test case #2256/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2257/2803" severity error;
    assert SOR = '0' report "Error in test case #2257/2803" severity error;
    assert SOL = '0' report "Error in test case #2257/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2258/2803" severity error;
    assert SOR = '0' report "Error in test case #2258/2803" severity error;
    assert SOL = '0' report "Error in test case #2258/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2259/2803" severity error;
    assert SOR = '0' report "Error in test case #2259/2803" severity error;
    assert SOL = '0' report "Error in test case #2259/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2260/2803" severity error;
    assert SOR = '0' report "Error in test case #2260/2803" severity error;
    assert SOL = '0' report "Error in test case #2260/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2261/2803" severity error;
    assert SOR = '0' report "Error in test case #2261/2803" severity error;
    assert SOL = '0' report "Error in test case #2261/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2262/2803" severity error;
    assert SOR = '0' report "Error in test case #2262/2803" severity error;
    assert SOL = '0' report "Error in test case #2262/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2263/2803" severity error;
    assert SOR = '0' report "Error in test case #2263/2803" severity error;
    assert SOL = '0' report "Error in test case #2263/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2264/2803" severity error;
    assert SOR = '0' report "Error in test case #2264/2803" severity error;
    assert SOL = '0' report "Error in test case #2264/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2265/2803" severity error;
    assert SOR = '0' report "Error in test case #2265/2803" severity error;
    assert SOL = '0' report "Error in test case #2265/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2266/2803" severity error;
    assert SOR = '0' report "Error in test case #2266/2803" severity error;
    assert SOL = '0' report "Error in test case #2266/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2267/2803" severity error;
    assert SOR = '0' report "Error in test case #2267/2803" severity error;
    assert SOL = '0' report "Error in test case #2267/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2268/2803" severity error;
    assert SOR = '0' report "Error in test case #2268/2803" severity error;
    assert SOL = '0' report "Error in test case #2268/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2269/2803" severity error;
    assert SOR = '0' report "Error in test case #2269/2803" severity error;
    assert SOL = '0' report "Error in test case #2269/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2270/2803" severity error;
    assert SOR = '0' report "Error in test case #2270/2803" severity error;
    assert SOL = '0' report "Error in test case #2270/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2271/2803" severity error;
    assert SOR = '0' report "Error in test case #2271/2803" severity error;
    assert SOL = '0' report "Error in test case #2271/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2272/2803" severity error;
    assert SOR = '0' report "Error in test case #2272/2803" severity error;
    assert SOL = '0' report "Error in test case #2272/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2273/2803" severity error;
    assert SOR = '0' report "Error in test case #2273/2803" severity error;
    assert SOL = '0' report "Error in test case #2273/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2274/2803" severity error;
    assert SOR = '0' report "Error in test case #2274/2803" severity error;
    assert SOL = '0' report "Error in test case #2274/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2275/2803" severity error;
    assert SOR = '0' report "Error in test case #2275/2803" severity error;
    assert SOL = '0' report "Error in test case #2275/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2276/2803" severity error;
    assert SOR = '0' report "Error in test case #2276/2803" severity error;
    assert SOL = '0' report "Error in test case #2276/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2277/2803" severity error;
    assert SOR = '0' report "Error in test case #2277/2803" severity error;
    assert SOL = '0' report "Error in test case #2277/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2278/2803" severity error;
    assert SOR = '0' report "Error in test case #2278/2803" severity error;
    assert SOL = '0' report "Error in test case #2278/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2279/2803" severity error;
    assert SOR = '0' report "Error in test case #2279/2803" severity error;
    assert SOL = '0' report "Error in test case #2279/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2280/2803" severity error;
    assert SOR = '0' report "Error in test case #2280/2803" severity error;
    assert SOL = '0' report "Error in test case #2280/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2281/2803" severity error;
    assert SOR = '0' report "Error in test case #2281/2803" severity error;
    assert SOL = '0' report "Error in test case #2281/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2282/2803" severity error;
    assert SOR = '0' report "Error in test case #2282/2803" severity error;
    assert SOL = '0' report "Error in test case #2282/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2283/2803" severity error;
    assert SOR = '0' report "Error in test case #2283/2803" severity error;
    assert SOL = '0' report "Error in test case #2283/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2284/2803" severity error;
    assert SOR = '0' report "Error in test case #2284/2803" severity error;
    assert SOL = '0' report "Error in test case #2284/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2285/2803" severity error;
    assert SOR = '0' report "Error in test case #2285/2803" severity error;
    assert SOL = '0' report "Error in test case #2285/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2286/2803" severity error;
    assert SOR = '0' report "Error in test case #2286/2803" severity error;
    assert SOL = '0' report "Error in test case #2286/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2287/2803" severity error;
    assert SOR = '0' report "Error in test case #2287/2803" severity error;
    assert SOL = '0' report "Error in test case #2287/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2288/2803" severity error;
    assert SOR = '0' report "Error in test case #2288/2803" severity error;
    assert SOL = '0' report "Error in test case #2288/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2289/2803" severity error;
    assert SOR = '0' report "Error in test case #2289/2803" severity error;
    assert SOL = '0' report "Error in test case #2289/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2290/2803" severity error;
    assert SOR = '0' report "Error in test case #2290/2803" severity error;
    assert SOL = '0' report "Error in test case #2290/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2291/2803" severity error;
    assert SOR = '0' report "Error in test case #2291/2803" severity error;
    assert SOL = '0' report "Error in test case #2291/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2292/2803" severity error;
    assert SOR = '0' report "Error in test case #2292/2803" severity error;
    assert SOL = '0' report "Error in test case #2292/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2293/2803" severity error;
    assert SOR = '0' report "Error in test case #2293/2803" severity error;
    assert SOL = '0' report "Error in test case #2293/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2294/2803" severity error;
    assert SOR = '0' report "Error in test case #2294/2803" severity error;
    assert SOL = '0' report "Error in test case #2294/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2295/2803" severity error;
    assert SOR = '0' report "Error in test case #2295/2803" severity error;
    assert SOL = '0' report "Error in test case #2295/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2296/2803" severity error;
    assert SOR = '0' report "Error in test case #2296/2803" severity error;
    assert SOL = '0' report "Error in test case #2296/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2297/2803" severity error;
    assert SOR = '0' report "Error in test case #2297/2803" severity error;
    assert SOL = '0' report "Error in test case #2297/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2298/2803" severity error;
    assert SOR = '0' report "Error in test case #2298/2803" severity error;
    assert SOL = '0' report "Error in test case #2298/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2299/2803" severity error;
    assert SOR = '0' report "Error in test case #2299/2803" severity error;
    assert SOL = '0' report "Error in test case #2299/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2300/2803" severity error;
    assert SOR = '0' report "Error in test case #2300/2803" severity error;
    assert SOL = '0' report "Error in test case #2300/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2301/2803" severity error;
    assert SOR = '0' report "Error in test case #2301/2803" severity error;
    assert SOL = '0' report "Error in test case #2301/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2302/2803" severity error;
    assert SOR = '0' report "Error in test case #2302/2803" severity error;
    assert SOL = '0' report "Error in test case #2302/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2303/2803" severity error;
    assert SOR = '0' report "Error in test case #2303/2803" severity error;
    assert SOL = '0' report "Error in test case #2303/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2304/2803" severity error;
    assert SOR = '0' report "Error in test case #2304/2803" severity error;
    assert SOL = '0' report "Error in test case #2304/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2305/2803" severity error;
    assert SOR = '0' report "Error in test case #2305/2803" severity error;
    assert SOL = '0' report "Error in test case #2305/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2306/2803" severity error;
    assert SOR = '0' report "Error in test case #2306/2803" severity error;
    assert SOL = '0' report "Error in test case #2306/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '0';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2307/2803" severity error;
    assert SOR = '0' report "Error in test case #2307/2803" severity error;
    assert SOL = '0' report "Error in test case #2307/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2308/2803" severity error;
    assert SOR = '0' report "Error in test case #2308/2803" severity error;
    assert SOL = '0' report "Error in test case #2308/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2309/2803" severity error;
    assert SOR = '0' report "Error in test case #2309/2803" severity error;
    assert SOL = '0' report "Error in test case #2309/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2310/2803" severity error;
    assert SOR = '0' report "Error in test case #2310/2803" severity error;
    assert SOL = '0' report "Error in test case #2310/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2311/2803" severity error;
    assert SOR = '0' report "Error in test case #2311/2803" severity error;
    assert SOL = '0' report "Error in test case #2311/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2312/2803" severity error;
    assert SOR = '0' report "Error in test case #2312/2803" severity error;
    assert SOL = '0' report "Error in test case #2312/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2313/2803" severity error;
    assert SOR = '0' report "Error in test case #2313/2803" severity error;
    assert SOL = '0' report "Error in test case #2313/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2314/2803" severity error;
    assert SOR = '0' report "Error in test case #2314/2803" severity error;
    assert SOL = '0' report "Error in test case #2314/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2315/2803" severity error;
    assert SOR = '0' report "Error in test case #2315/2803" severity error;
    assert SOL = '0' report "Error in test case #2315/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2316/2803" severity error;
    assert SOR = '0' report "Error in test case #2316/2803" severity error;
    assert SOL = '0' report "Error in test case #2316/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2317/2803" severity error;
    assert SOR = '0' report "Error in test case #2317/2803" severity error;
    assert SOL = '0' report "Error in test case #2317/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2318/2803" severity error;
    assert SOR = '0' report "Error in test case #2318/2803" severity error;
    assert SOL = '0' report "Error in test case #2318/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2319/2803" severity error;
    assert SOR = '0' report "Error in test case #2319/2803" severity error;
    assert SOL = '0' report "Error in test case #2319/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2320/2803" severity error;
    assert SOR = '0' report "Error in test case #2320/2803" severity error;
    assert SOL = '0' report "Error in test case #2320/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2321/2803" severity error;
    assert SOR = '0' report "Error in test case #2321/2803" severity error;
    assert SOL = '0' report "Error in test case #2321/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2322/2803" severity error;
    assert SOR = '0' report "Error in test case #2322/2803" severity error;
    assert SOL = '0' report "Error in test case #2322/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2323/2803" severity error;
    assert SOR = '0' report "Error in test case #2323/2803" severity error;
    assert SOL = '0' report "Error in test case #2323/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2324/2803" severity error;
    assert SOR = '0' report "Error in test case #2324/2803" severity error;
    assert SOL = '0' report "Error in test case #2324/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2325/2803" severity error;
    assert SOR = '0' report "Error in test case #2325/2803" severity error;
    assert SOL = '0' report "Error in test case #2325/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2326/2803" severity error;
    assert SOR = '0' report "Error in test case #2326/2803" severity error;
    assert SOL = '0' report "Error in test case #2326/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2327/2803" severity error;
    assert SOR = '0' report "Error in test case #2327/2803" severity error;
    assert SOL = '0' report "Error in test case #2327/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2328/2803" severity error;
    assert SOR = '0' report "Error in test case #2328/2803" severity error;
    assert SOL = '0' report "Error in test case #2328/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2329/2803" severity error;
    assert SOR = '0' report "Error in test case #2329/2803" severity error;
    assert SOL = '0' report "Error in test case #2329/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2330/2803" severity error;
    assert SOR = '0' report "Error in test case #2330/2803" severity error;
    assert SOL = '0' report "Error in test case #2330/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2331/2803" severity error;
    assert SOR = '0' report "Error in test case #2331/2803" severity error;
    assert SOL = '0' report "Error in test case #2331/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2332/2803" severity error;
    assert SOR = '0' report "Error in test case #2332/2803" severity error;
    assert SOL = '0' report "Error in test case #2332/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2333/2803" severity error;
    assert SOR = '0' report "Error in test case #2333/2803" severity error;
    assert SOL = '0' report "Error in test case #2333/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2334/2803" severity error;
    assert SOR = '0' report "Error in test case #2334/2803" severity error;
    assert SOL = '0' report "Error in test case #2334/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2335/2803" severity error;
    assert SOR = '0' report "Error in test case #2335/2803" severity error;
    assert SOL = '0' report "Error in test case #2335/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2336/2803" severity error;
    assert SOR = '0' report "Error in test case #2336/2803" severity error;
    assert SOL = '0' report "Error in test case #2336/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2337/2803" severity error;
    assert SOR = '0' report "Error in test case #2337/2803" severity error;
    assert SOL = '0' report "Error in test case #2337/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2338/2803" severity error;
    assert SOR = '0' report "Error in test case #2338/2803" severity error;
    assert SOL = '0' report "Error in test case #2338/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2339/2803" severity error;
    assert SOR = '0' report "Error in test case #2339/2803" severity error;
    assert SOL = '0' report "Error in test case #2339/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2340/2803" severity error;
    assert SOR = '0' report "Error in test case #2340/2803" severity error;
    assert SOL = '0' report "Error in test case #2340/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2341/2803" severity error;
    assert SOR = '0' report "Error in test case #2341/2803" severity error;
    assert SOL = '0' report "Error in test case #2341/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2342/2803" severity error;
    assert SOR = '0' report "Error in test case #2342/2803" severity error;
    assert SOL = '0' report "Error in test case #2342/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2343/2803" severity error;
    assert SOR = '0' report "Error in test case #2343/2803" severity error;
    assert SOL = '0' report "Error in test case #2343/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2344/2803" severity error;
    assert SOR = '0' report "Error in test case #2344/2803" severity error;
    assert SOL = '0' report "Error in test case #2344/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2345/2803" severity error;
    assert SOR = '0' report "Error in test case #2345/2803" severity error;
    assert SOL = '0' report "Error in test case #2345/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2346/2803" severity error;
    assert SOR = '0' report "Error in test case #2346/2803" severity error;
    assert SOL = '0' report "Error in test case #2346/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2347/2803" severity error;
    assert SOR = '0' report "Error in test case #2347/2803" severity error;
    assert SOL = '0' report "Error in test case #2347/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2348/2803" severity error;
    assert SOR = '0' report "Error in test case #2348/2803" severity error;
    assert SOL = '0' report "Error in test case #2348/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2349/2803" severity error;
    assert SOR = '0' report "Error in test case #2349/2803" severity error;
    assert SOL = '0' report "Error in test case #2349/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2350/2803" severity error;
    assert SOR = '0' report "Error in test case #2350/2803" severity error;
    assert SOL = '0' report "Error in test case #2350/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2351/2803" severity error;
    assert SOR = '0' report "Error in test case #2351/2803" severity error;
    assert SOL = '0' report "Error in test case #2351/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2352/2803" severity error;
    assert SOR = '0' report "Error in test case #2352/2803" severity error;
    assert SOL = '0' report "Error in test case #2352/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2353/2803" severity error;
    assert SOR = '0' report "Error in test case #2353/2803" severity error;
    assert SOL = '0' report "Error in test case #2353/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2354/2803" severity error;
    assert SOR = '0' report "Error in test case #2354/2803" severity error;
    assert SOL = '0' report "Error in test case #2354/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2355/2803" severity error;
    assert SOR = '0' report "Error in test case #2355/2803" severity error;
    assert SOL = '0' report "Error in test case #2355/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2356/2803" severity error;
    assert SOR = '0' report "Error in test case #2356/2803" severity error;
    assert SOL = '0' report "Error in test case #2356/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2357/2803" severity error;
    assert SOR = '0' report "Error in test case #2357/2803" severity error;
    assert SOL = '0' report "Error in test case #2357/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2358/2803" severity error;
    assert SOR = '0' report "Error in test case #2358/2803" severity error;
    assert SOL = '0' report "Error in test case #2358/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2359/2803" severity error;
    assert SOR = '0' report "Error in test case #2359/2803" severity error;
    assert SOL = '0' report "Error in test case #2359/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2360/2803" severity error;
    assert SOR = '0' report "Error in test case #2360/2803" severity error;
    assert SOL = '0' report "Error in test case #2360/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2361/2803" severity error;
    assert SOR = '0' report "Error in test case #2361/2803" severity error;
    assert SOL = '0' report "Error in test case #2361/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2362/2803" severity error;
    assert SOR = '0' report "Error in test case #2362/2803" severity error;
    assert SOL = '0' report "Error in test case #2362/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2363/2803" severity error;
    assert SOR = '0' report "Error in test case #2363/2803" severity error;
    assert SOL = '0' report "Error in test case #2363/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2364/2803" severity error;
    assert SOR = '0' report "Error in test case #2364/2803" severity error;
    assert SOL = '0' report "Error in test case #2364/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2365/2803" severity error;
    assert SOR = '0' report "Error in test case #2365/2803" severity error;
    assert SOL = '0' report "Error in test case #2365/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2366/2803" severity error;
    assert SOR = '0' report "Error in test case #2366/2803" severity error;
    assert SOL = '0' report "Error in test case #2366/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2367/2803" severity error;
    assert SOR = '0' report "Error in test case #2367/2803" severity error;
    assert SOL = '0' report "Error in test case #2367/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2368/2803" severity error;
    assert SOR = '0' report "Error in test case #2368/2803" severity error;
    assert SOL = '0' report "Error in test case #2368/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2369/2803" severity error;
    assert SOR = '0' report "Error in test case #2369/2803" severity error;
    assert SOL = '0' report "Error in test case #2369/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2370/2803" severity error;
    assert SOR = '0' report "Error in test case #2370/2803" severity error;
    assert SOL = '0' report "Error in test case #2370/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2371/2803" severity error;
    assert SOR = '0' report "Error in test case #2371/2803" severity error;
    assert SOL = '0' report "Error in test case #2371/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2372/2803" severity error;
    assert SOR = '0' report "Error in test case #2372/2803" severity error;
    assert SOL = '0' report "Error in test case #2372/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2373/2803" severity error;
    assert SOR = '0' report "Error in test case #2373/2803" severity error;
    assert SOL = '0' report "Error in test case #2373/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2374/2803" severity error;
    assert SOR = '0' report "Error in test case #2374/2803" severity error;
    assert SOL = '0' report "Error in test case #2374/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2375/2803" severity error;
    assert SOR = '0' report "Error in test case #2375/2803" severity error;
    assert SOL = '0' report "Error in test case #2375/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2376/2803" severity error;
    assert SOR = '0' report "Error in test case #2376/2803" severity error;
    assert SOL = '0' report "Error in test case #2376/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2377/2803" severity error;
    assert SOR = '0' report "Error in test case #2377/2803" severity error;
    assert SOL = '0' report "Error in test case #2377/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2378/2803" severity error;
    assert SOR = '0' report "Error in test case #2378/2803" severity error;
    assert SOL = '0' report "Error in test case #2378/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2379/2803" severity error;
    assert SOR = '0' report "Error in test case #2379/2803" severity error;
    assert SOL = '0' report "Error in test case #2379/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2380/2803" severity error;
    assert SOR = '0' report "Error in test case #2380/2803" severity error;
    assert SOL = '0' report "Error in test case #2380/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2381/2803" severity error;
    assert SOR = '0' report "Error in test case #2381/2803" severity error;
    assert SOL = '0' report "Error in test case #2381/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2382/2803" severity error;
    assert SOR = '0' report "Error in test case #2382/2803" severity error;
    assert SOL = '0' report "Error in test case #2382/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2383/2803" severity error;
    assert SOR = '0' report "Error in test case #2383/2803" severity error;
    assert SOL = '0' report "Error in test case #2383/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2384/2803" severity error;
    assert SOR = '0' report "Error in test case #2384/2803" severity error;
    assert SOL = '0' report "Error in test case #2384/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2385/2803" severity error;
    assert SOR = '0' report "Error in test case #2385/2803" severity error;
    assert SOL = '0' report "Error in test case #2385/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2386/2803" severity error;
    assert SOR = '0' report "Error in test case #2386/2803" severity error;
    assert SOL = '0' report "Error in test case #2386/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2387/2803" severity error;
    assert SOR = '0' report "Error in test case #2387/2803" severity error;
    assert SOL = '0' report "Error in test case #2387/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2388/2803" severity error;
    assert SOR = '0' report "Error in test case #2388/2803" severity error;
    assert SOL = '0' report "Error in test case #2388/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2389/2803" severity error;
    assert SOR = '0' report "Error in test case #2389/2803" severity error;
    assert SOL = '0' report "Error in test case #2389/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2390/2803" severity error;
    assert SOR = '0' report "Error in test case #2390/2803" severity error;
    assert SOL = '0' report "Error in test case #2390/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2391/2803" severity error;
    assert SOR = '0' report "Error in test case #2391/2803" severity error;
    assert SOL = '0' report "Error in test case #2391/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2392/2803" severity error;
    assert SOR = '0' report "Error in test case #2392/2803" severity error;
    assert SOL = '0' report "Error in test case #2392/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2393/2803" severity error;
    assert SOR = '0' report "Error in test case #2393/2803" severity error;
    assert SOL = '0' report "Error in test case #2393/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2394/2803" severity error;
    assert SOR = '0' report "Error in test case #2394/2803" severity error;
    assert SOL = '0' report "Error in test case #2394/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2395/2803" severity error;
    assert SOR = '0' report "Error in test case #2395/2803" severity error;
    assert SOL = '0' report "Error in test case #2395/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2396/2803" severity error;
    assert SOR = '0' report "Error in test case #2396/2803" severity error;
    assert SOL = '0' report "Error in test case #2396/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2397/2803" severity error;
    assert SOR = '0' report "Error in test case #2397/2803" severity error;
    assert SOL = '0' report "Error in test case #2397/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2398/2803" severity error;
    assert SOR = '0' report "Error in test case #2398/2803" severity error;
    assert SOL = '0' report "Error in test case #2398/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2399/2803" severity error;
    assert SOR = '0' report "Error in test case #2399/2803" severity error;
    assert SOL = '0' report "Error in test case #2399/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2400/2803" severity error;
    assert SOR = '1' report "Error in test case #2400/2803" severity error;
    assert SOL = '1' report "Error in test case #2400/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2401/2803" severity error;
    assert SOR = '1' report "Error in test case #2401/2803" severity error;
    assert SOL = '1' report "Error in test case #2401/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2402/2803" severity error;
    assert SOR = '1' report "Error in test case #2402/2803" severity error;
    assert SOL = '1' report "Error in test case #2402/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "101";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2403/2803" severity error;
    assert SOR = '1' report "Error in test case #2403/2803" severity error;
    assert SOL = '1' report "Error in test case #2403/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2404/2803" severity error;
    assert SOR = '1' report "Error in test case #2404/2803" severity error;
    assert SOL = '1' report "Error in test case #2404/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2405/2803" severity error;
    assert SOR = '1' report "Error in test case #2405/2803" severity error;
    assert SOL = '1' report "Error in test case #2405/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2406/2803" severity error;
    assert SOR = '1' report "Error in test case #2406/2803" severity error;
    assert SOL = '1' report "Error in test case #2406/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2407/2803" severity error;
    assert SOR = '1' report "Error in test case #2407/2803" severity error;
    assert SOL = '1' report "Error in test case #2407/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2408/2803" severity error;
    assert SOR = '1' report "Error in test case #2408/2803" severity error;
    assert SOL = '1' report "Error in test case #2408/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2409/2803" severity error;
    assert SOR = '1' report "Error in test case #2409/2803" severity error;
    assert SOL = '1' report "Error in test case #2409/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2410/2803" severity error;
    assert SOR = '1' report "Error in test case #2410/2803" severity error;
    assert SOL = '1' report "Error in test case #2410/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2411/2803" severity error;
    assert SOR = '1' report "Error in test case #2411/2803" severity error;
    assert SOL = '1' report "Error in test case #2411/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2412/2803" severity error;
    assert SOR = '1' report "Error in test case #2412/2803" severity error;
    assert SOL = '1' report "Error in test case #2412/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2413/2803" severity error;
    assert SOR = '1' report "Error in test case #2413/2803" severity error;
    assert SOL = '1' report "Error in test case #2413/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2414/2803" severity error;
    assert SOR = '1' report "Error in test case #2414/2803" severity error;
    assert SOL = '1' report "Error in test case #2414/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2415/2803" severity error;
    assert SOR = '1' report "Error in test case #2415/2803" severity error;
    assert SOL = '1' report "Error in test case #2415/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2416/2803" severity error;
    assert SOR = '1' report "Error in test case #2416/2803" severity error;
    assert SOL = '1' report "Error in test case #2416/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2417/2803" severity error;
    assert SOR = '1' report "Error in test case #2417/2803" severity error;
    assert SOL = '1' report "Error in test case #2417/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2418/2803" severity error;
    assert SOR = '1' report "Error in test case #2418/2803" severity error;
    assert SOL = '1' report "Error in test case #2418/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2419/2803" severity error;
    assert SOR = '1' report "Error in test case #2419/2803" severity error;
    assert SOL = '1' report "Error in test case #2419/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2420/2803" severity error;
    assert SOR = '1' report "Error in test case #2420/2803" severity error;
    assert SOL = '1' report "Error in test case #2420/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2421/2803" severity error;
    assert SOR = '1' report "Error in test case #2421/2803" severity error;
    assert SOL = '1' report "Error in test case #2421/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2422/2803" severity error;
    assert SOR = '0' report "Error in test case #2422/2803" severity error;
    assert SOL = '0' report "Error in test case #2422/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2423/2803" severity error;
    assert SOR = '0' report "Error in test case #2423/2803" severity error;
    assert SOL = '0' report "Error in test case #2423/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2424/2803" severity error;
    assert SOR = '0' report "Error in test case #2424/2803" severity error;
    assert SOL = '0' report "Error in test case #2424/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2425/2803" severity error;
    assert SOR = '0' report "Error in test case #2425/2803" severity error;
    assert SOL = '0' report "Error in test case #2425/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2426/2803" severity error;
    assert SOR = '0' report "Error in test case #2426/2803" severity error;
    assert SOL = '0' report "Error in test case #2426/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2427/2803" severity error;
    assert SOR = '0' report "Error in test case #2427/2803" severity error;
    assert SOL = '0' report "Error in test case #2427/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2428/2803" severity error;
    assert SOR = '0' report "Error in test case #2428/2803" severity error;
    assert SOL = '0' report "Error in test case #2428/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2429/2803" severity error;
    assert SOR = '0' report "Error in test case #2429/2803" severity error;
    assert SOL = '0' report "Error in test case #2429/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2430/2803" severity error;
    assert SOR = '0' report "Error in test case #2430/2803" severity error;
    assert SOL = '0' report "Error in test case #2430/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2431/2803" severity error;
    assert SOR = '0' report "Error in test case #2431/2803" severity error;
    assert SOL = '0' report "Error in test case #2431/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2432/2803" severity error;
    assert SOR = '0' report "Error in test case #2432/2803" severity error;
    assert SOL = '0' report "Error in test case #2432/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2433/2803" severity error;
    assert SOR = '0' report "Error in test case #2433/2803" severity error;
    assert SOL = '0' report "Error in test case #2433/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2434/2803" severity error;
    assert SOR = '0' report "Error in test case #2434/2803" severity error;
    assert SOL = '0' report "Error in test case #2434/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2435/2803" severity error;
    assert SOR = '0' report "Error in test case #2435/2803" severity error;
    assert SOL = '0' report "Error in test case #2435/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2436/2803" severity error;
    assert SOR = '0' report "Error in test case #2436/2803" severity error;
    assert SOL = '0' report "Error in test case #2436/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2437/2803" severity error;
    assert SOR = '0' report "Error in test case #2437/2803" severity error;
    assert SOL = '0' report "Error in test case #2437/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2438/2803" severity error;
    assert SOR = '0' report "Error in test case #2438/2803" severity error;
    assert SOL = '0' report "Error in test case #2438/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2439/2803" severity error;
    assert SOR = '0' report "Error in test case #2439/2803" severity error;
    assert SOL = '0' report "Error in test case #2439/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2440/2803" severity error;
    assert SOR = '0' report "Error in test case #2440/2803" severity error;
    assert SOL = '0' report "Error in test case #2440/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2441/2803" severity error;
    assert SOR = '0' report "Error in test case #2441/2803" severity error;
    assert SOL = '0' report "Error in test case #2441/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2442/2803" severity error;
    assert SOR = '0' report "Error in test case #2442/2803" severity error;
    assert SOL = '0' report "Error in test case #2442/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2443/2803" severity error;
    assert SOR = '0' report "Error in test case #2443/2803" severity error;
    assert SOL = '0' report "Error in test case #2443/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2444/2803" severity error;
    assert SOR = '0' report "Error in test case #2444/2803" severity error;
    assert SOL = '0' report "Error in test case #2444/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2445/2803" severity error;
    assert SOR = '0' report "Error in test case #2445/2803" severity error;
    assert SOL = '0' report "Error in test case #2445/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2446/2803" severity error;
    assert SOR = '1' report "Error in test case #2446/2803" severity error;
    assert SOL = '1' report "Error in test case #2446/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2447/2803" severity error;
    assert SOR = '1' report "Error in test case #2447/2803" severity error;
    assert SOL = '1' report "Error in test case #2447/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2448/2803" severity error;
    assert SOR = '1' report "Error in test case #2448/2803" severity error;
    assert SOL = '1' report "Error in test case #2448/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2449/2803" severity error;
    assert SOR = '1' report "Error in test case #2449/2803" severity error;
    assert SOL = '1' report "Error in test case #2449/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2450/2803" severity error;
    assert SOR = '1' report "Error in test case #2450/2803" severity error;
    assert SOL = '1' report "Error in test case #2450/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2451/2803" severity error;
    assert SOR = '1' report "Error in test case #2451/2803" severity error;
    assert SOL = '1' report "Error in test case #2451/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2452/2803" severity error;
    assert SOR = '1' report "Error in test case #2452/2803" severity error;
    assert SOL = '1' report "Error in test case #2452/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2453/2803" severity error;
    assert SOR = '1' report "Error in test case #2453/2803" severity error;
    assert SOL = '1' report "Error in test case #2453/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2454/2803" severity error;
    assert SOR = '1' report "Error in test case #2454/2803" severity error;
    assert SOL = '1' report "Error in test case #2454/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2455/2803" severity error;
    assert SOR = '1' report "Error in test case #2455/2803" severity error;
    assert SOL = '1' report "Error in test case #2455/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2456/2803" severity error;
    assert SOR = '1' report "Error in test case #2456/2803" severity error;
    assert SOL = '1' report "Error in test case #2456/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2457/2803" severity error;
    assert SOR = '1' report "Error in test case #2457/2803" severity error;
    assert SOL = '1' report "Error in test case #2457/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2458/2803" severity error;
    assert SOR = '1' report "Error in test case #2458/2803" severity error;
    assert SOL = '1' report "Error in test case #2458/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2459/2803" severity error;
    assert SOR = '1' report "Error in test case #2459/2803" severity error;
    assert SOL = '1' report "Error in test case #2459/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2460/2803" severity error;
    assert SOR = '1' report "Error in test case #2460/2803" severity error;
    assert SOL = '1' report "Error in test case #2460/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2461/2803" severity error;
    assert SOR = '1' report "Error in test case #2461/2803" severity error;
    assert SOL = '1' report "Error in test case #2461/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2462/2803" severity error;
    assert SOR = '1' report "Error in test case #2462/2803" severity error;
    assert SOL = '1' report "Error in test case #2462/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2463/2803" severity error;
    assert SOR = '1' report "Error in test case #2463/2803" severity error;
    assert SOL = '1' report "Error in test case #2463/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2464/2803" severity error;
    assert SOR = '1' report "Error in test case #2464/2803" severity error;
    assert SOL = '1' report "Error in test case #2464/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2465/2803" severity error;
    assert SOR = '1' report "Error in test case #2465/2803" severity error;
    assert SOL = '1' report "Error in test case #2465/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2466/2803" severity error;
    assert SOR = '1' report "Error in test case #2466/2803" severity error;
    assert SOL = '1' report "Error in test case #2466/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2467/2803" severity error;
    assert SOR = '1' report "Error in test case #2467/2803" severity error;
    assert SOL = '1' report "Error in test case #2467/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2468/2803" severity error;
    assert SOR = '1' report "Error in test case #2468/2803" severity error;
    assert SOL = '1' report "Error in test case #2468/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2469/2803" severity error;
    assert SOR = '1' report "Error in test case #2469/2803" severity error;
    assert SOL = '1' report "Error in test case #2469/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2470/2803" severity error;
    assert SOR = '1' report "Error in test case #2470/2803" severity error;
    assert SOL = '1' report "Error in test case #2470/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2471/2803" severity error;
    assert SOR = '1' report "Error in test case #2471/2803" severity error;
    assert SOL = '1' report "Error in test case #2471/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2472/2803" severity error;
    assert SOR = '1' report "Error in test case #2472/2803" severity error;
    assert SOL = '1' report "Error in test case #2472/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2473/2803" severity error;
    assert SOR = '1' report "Error in test case #2473/2803" severity error;
    assert SOL = '1' report "Error in test case #2473/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2474/2803" severity error;
    assert SOR = '1' report "Error in test case #2474/2803" severity error;
    assert SOL = '1' report "Error in test case #2474/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2475/2803" severity error;
    assert SOR = '1' report "Error in test case #2475/2803" severity error;
    assert SOL = '1' report "Error in test case #2475/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2476/2803" severity error;
    assert SOR = '1' report "Error in test case #2476/2803" severity error;
    assert SOL = '1' report "Error in test case #2476/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2477/2803" severity error;
    assert SOR = '1' report "Error in test case #2477/2803" severity error;
    assert SOL = '1' report "Error in test case #2477/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2478/2803" severity error;
    assert SOR = '1' report "Error in test case #2478/2803" severity error;
    assert SOL = '1' report "Error in test case #2478/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2479/2803" severity error;
    assert SOR = '1' report "Error in test case #2479/2803" severity error;
    assert SOL = '1' report "Error in test case #2479/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2480/2803" severity error;
    assert SOR = '1' report "Error in test case #2480/2803" severity error;
    assert SOL = '1' report "Error in test case #2480/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2481/2803" severity error;
    assert SOR = '1' report "Error in test case #2481/2803" severity error;
    assert SOL = '1' report "Error in test case #2481/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2482/2803" severity error;
    assert SOR = '1' report "Error in test case #2482/2803" severity error;
    assert SOL = '1' report "Error in test case #2482/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2483/2803" severity error;
    assert SOR = '1' report "Error in test case #2483/2803" severity error;
    assert SOL = '1' report "Error in test case #2483/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2484/2803" severity error;
    assert SOR = '1' report "Error in test case #2484/2803" severity error;
    assert SOL = '1' report "Error in test case #2484/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2485/2803" severity error;
    assert SOR = '1' report "Error in test case #2485/2803" severity error;
    assert SOL = '1' report "Error in test case #2485/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2486/2803" severity error;
    assert SOR = '0' report "Error in test case #2486/2803" severity error;
    assert SOL = '0' report "Error in test case #2486/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2487/2803" severity error;
    assert SOR = '0' report "Error in test case #2487/2803" severity error;
    assert SOL = '0' report "Error in test case #2487/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2488/2803" severity error;
    assert SOR = '0' report "Error in test case #2488/2803" severity error;
    assert SOL = '0' report "Error in test case #2488/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2489/2803" severity error;
    assert SOR = '0' report "Error in test case #2489/2803" severity error;
    assert SOL = '0' report "Error in test case #2489/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2490/2803" severity error;
    assert SOR = '0' report "Error in test case #2490/2803" severity error;
    assert SOL = '0' report "Error in test case #2490/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2491/2803" severity error;
    assert SOR = '0' report "Error in test case #2491/2803" severity error;
    assert SOL = '0' report "Error in test case #2491/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2492/2803" severity error;
    assert SOR = '0' report "Error in test case #2492/2803" severity error;
    assert SOL = '0' report "Error in test case #2492/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2493/2803" severity error;
    assert SOR = '0' report "Error in test case #2493/2803" severity error;
    assert SOL = '0' report "Error in test case #2493/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2494/2803" severity error;
    assert SOR = '0' report "Error in test case #2494/2803" severity error;
    assert SOL = '0' report "Error in test case #2494/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2495/2803" severity error;
    assert SOR = '0' report "Error in test case #2495/2803" severity error;
    assert SOL = '0' report "Error in test case #2495/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2496/2803" severity error;
    assert SOR = '0' report "Error in test case #2496/2803" severity error;
    assert SOL = '0' report "Error in test case #2496/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2497/2803" severity error;
    assert SOR = '0' report "Error in test case #2497/2803" severity error;
    assert SOL = '0' report "Error in test case #2497/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2498/2803" severity error;
    assert SOR = '0' report "Error in test case #2498/2803" severity error;
    assert SOL = '0' report "Error in test case #2498/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2499/2803" severity error;
    assert SOR = '0' report "Error in test case #2499/2803" severity error;
    assert SOL = '0' report "Error in test case #2499/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2500/2803" severity error;
    assert SOR = '0' report "Error in test case #2500/2803" severity error;
    assert SOL = '0' report "Error in test case #2500/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2501/2803" severity error;
    assert SOR = '0' report "Error in test case #2501/2803" severity error;
    assert SOL = '0' report "Error in test case #2501/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2502/2803" severity error;
    assert SOR = '0' report "Error in test case #2502/2803" severity error;
    assert SOL = '0' report "Error in test case #2502/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2503/2803" severity error;
    assert SOR = '0' report "Error in test case #2503/2803" severity error;
    assert SOL = '0' report "Error in test case #2503/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2504/2803" severity error;
    assert SOR = '0' report "Error in test case #2504/2803" severity error;
    assert SOL = '0' report "Error in test case #2504/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2505/2803" severity error;
    assert SOR = '0' report "Error in test case #2505/2803" severity error;
    assert SOL = '0' report "Error in test case #2505/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2506/2803" severity error;
    assert SOR = '0' report "Error in test case #2506/2803" severity error;
    assert SOL = '0' report "Error in test case #2506/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2507/2803" severity error;
    assert SOR = '0' report "Error in test case #2507/2803" severity error;
    assert SOL = '0' report "Error in test case #2507/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2508/2803" severity error;
    assert SOR = '0' report "Error in test case #2508/2803" severity error;
    assert SOL = '0' report "Error in test case #2508/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2509/2803" severity error;
    assert SOR = '0' report "Error in test case #2509/2803" severity error;
    assert SOL = '0' report "Error in test case #2509/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2510/2803" severity error;
    assert SOR = '1' report "Error in test case #2510/2803" severity error;
    assert SOL = '1' report "Error in test case #2510/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2511/2803" severity error;
    assert SOR = '1' report "Error in test case #2511/2803" severity error;
    assert SOL = '1' report "Error in test case #2511/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2512/2803" severity error;
    assert SOR = '1' report "Error in test case #2512/2803" severity error;
    assert SOL = '1' report "Error in test case #2512/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2513/2803" severity error;
    assert SOR = '1' report "Error in test case #2513/2803" severity error;
    assert SOL = '1' report "Error in test case #2513/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2514/2803" severity error;
    assert SOR = '1' report "Error in test case #2514/2803" severity error;
    assert SOL = '1' report "Error in test case #2514/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2515/2803" severity error;
    assert SOR = '1' report "Error in test case #2515/2803" severity error;
    assert SOL = '1' report "Error in test case #2515/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2516/2803" severity error;
    assert SOR = '1' report "Error in test case #2516/2803" severity error;
    assert SOL = '1' report "Error in test case #2516/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2517/2803" severity error;
    assert SOR = '1' report "Error in test case #2517/2803" severity error;
    assert SOL = '1' report "Error in test case #2517/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2518/2803" severity error;
    assert SOR = '1' report "Error in test case #2518/2803" severity error;
    assert SOL = '1' report "Error in test case #2518/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2519/2803" severity error;
    assert SOR = '1' report "Error in test case #2519/2803" severity error;
    assert SOL = '1' report "Error in test case #2519/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2520/2803" severity error;
    assert SOR = '1' report "Error in test case #2520/2803" severity error;
    assert SOL = '1' report "Error in test case #2520/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2521/2803" severity error;
    assert SOR = '1' report "Error in test case #2521/2803" severity error;
    assert SOL = '1' report "Error in test case #2521/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2522/2803" severity error;
    assert SOR = '1' report "Error in test case #2522/2803" severity error;
    assert SOL = '1' report "Error in test case #2522/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2523/2803" severity error;
    assert SOR = '1' report "Error in test case #2523/2803" severity error;
    assert SOL = '1' report "Error in test case #2523/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2524/2803" severity error;
    assert SOR = '1' report "Error in test case #2524/2803" severity error;
    assert SOL = '1' report "Error in test case #2524/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2525/2803" severity error;
    assert SOR = '1' report "Error in test case #2525/2803" severity error;
    assert SOL = '1' report "Error in test case #2525/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2526/2803" severity error;
    assert SOR = '1' report "Error in test case #2526/2803" severity error;
    assert SOL = '1' report "Error in test case #2526/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2527/2803" severity error;
    assert SOR = '1' report "Error in test case #2527/2803" severity error;
    assert SOL = '1' report "Error in test case #2527/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2528/2803" severity error;
    assert SOR = '1' report "Error in test case #2528/2803" severity error;
    assert SOL = '1' report "Error in test case #2528/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2529/2803" severity error;
    assert SOR = '1' report "Error in test case #2529/2803" severity error;
    assert SOL = '1' report "Error in test case #2529/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2530/2803" severity error;
    assert SOR = '1' report "Error in test case #2530/2803" severity error;
    assert SOL = '1' report "Error in test case #2530/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2531/2803" severity error;
    assert SOR = '1' report "Error in test case #2531/2803" severity error;
    assert SOL = '1' report "Error in test case #2531/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2532/2803" severity error;
    assert SOR = '1' report "Error in test case #2532/2803" severity error;
    assert SOL = '1' report "Error in test case #2532/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2533/2803" severity error;
    assert SOR = '1' report "Error in test case #2533/2803" severity error;
    assert SOL = '1' report "Error in test case #2533/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2534/2803" severity error;
    assert SOR = '1' report "Error in test case #2534/2803" severity error;
    assert SOL = '1' report "Error in test case #2534/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2535/2803" severity error;
    assert SOR = '1' report "Error in test case #2535/2803" severity error;
    assert SOL = '1' report "Error in test case #2535/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2536/2803" severity error;
    assert SOR = '1' report "Error in test case #2536/2803" severity error;
    assert SOL = '1' report "Error in test case #2536/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2537/2803" severity error;
    assert SOR = '1' report "Error in test case #2537/2803" severity error;
    assert SOL = '1' report "Error in test case #2537/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2538/2803" severity error;
    assert SOR = '1' report "Error in test case #2538/2803" severity error;
    assert SOL = '1' report "Error in test case #2538/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2539/2803" severity error;
    assert SOR = '1' report "Error in test case #2539/2803" severity error;
    assert SOL = '1' report "Error in test case #2539/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2540/2803" severity error;
    assert SOR = '1' report "Error in test case #2540/2803" severity error;
    assert SOL = '1' report "Error in test case #2540/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2541/2803" severity error;
    assert SOR = '1' report "Error in test case #2541/2803" severity error;
    assert SOL = '1' report "Error in test case #2541/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2542/2803" severity error;
    assert SOR = '1' report "Error in test case #2542/2803" severity error;
    assert SOL = '1' report "Error in test case #2542/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2543/2803" severity error;
    assert SOR = '1' report "Error in test case #2543/2803" severity error;
    assert SOL = '1' report "Error in test case #2543/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2544/2803" severity error;
    assert SOR = '1' report "Error in test case #2544/2803" severity error;
    assert SOL = '1' report "Error in test case #2544/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2545/2803" severity error;
    assert SOR = '1' report "Error in test case #2545/2803" severity error;
    assert SOL = '1' report "Error in test case #2545/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2546/2803" severity error;
    assert SOR = '1' report "Error in test case #2546/2803" severity error;
    assert SOL = '1' report "Error in test case #2546/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2547/2803" severity error;
    assert SOR = '1' report "Error in test case #2547/2803" severity error;
    assert SOL = '1' report "Error in test case #2547/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2548/2803" severity error;
    assert SOR = '1' report "Error in test case #2548/2803" severity error;
    assert SOL = '1' report "Error in test case #2548/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2549/2803" severity error;
    assert SOR = '1' report "Error in test case #2549/2803" severity error;
    assert SOL = '1' report "Error in test case #2549/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2550/2803" severity error;
    assert SOR = '1' report "Error in test case #2550/2803" severity error;
    assert SOL = '1' report "Error in test case #2550/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2551/2803" severity error;
    assert SOR = '1' report "Error in test case #2551/2803" severity error;
    assert SOL = '1' report "Error in test case #2551/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2552/2803" severity error;
    assert SOR = '1' report "Error in test case #2552/2803" severity error;
    assert SOL = '1' report "Error in test case #2552/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2553/2803" severity error;
    assert SOR = '1' report "Error in test case #2553/2803" severity error;
    assert SOL = '1' report "Error in test case #2553/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2554/2803" severity error;
    assert SOR = '1' report "Error in test case #2554/2803" severity error;
    assert SOL = '1' report "Error in test case #2554/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2555/2803" severity error;
    assert SOR = '1' report "Error in test case #2555/2803" severity error;
    assert SOL = '1' report "Error in test case #2555/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2556/2803" severity error;
    assert SOR = '1' report "Error in test case #2556/2803" severity error;
    assert SOL = '1' report "Error in test case #2556/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2557/2803" severity error;
    assert SOR = '1' report "Error in test case #2557/2803" severity error;
    assert SOL = '1' report "Error in test case #2557/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2558/2803" severity error;
    assert SOR = '1' report "Error in test case #2558/2803" severity error;
    assert SOL = '1' report "Error in test case #2558/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2559/2803" severity error;
    assert SOR = '1' report "Error in test case #2559/2803" severity error;
    assert SOL = '1' report "Error in test case #2559/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2560/2803" severity error;
    assert SOR = '1' report "Error in test case #2560/2803" severity error;
    assert SOL = '1' report "Error in test case #2560/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2561/2803" severity error;
    assert SOR = '1' report "Error in test case #2561/2803" severity error;
    assert SOL = '1' report "Error in test case #2561/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2562/2803" severity error;
    assert SOR = '1' report "Error in test case #2562/2803" severity error;
    assert SOL = '1' report "Error in test case #2562/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2563/2803" severity error;
    assert SOR = '1' report "Error in test case #2563/2803" severity error;
    assert SOL = '1' report "Error in test case #2563/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2564/2803" severity error;
    assert SOR = '1' report "Error in test case #2564/2803" severity error;
    assert SOL = '1' report "Error in test case #2564/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2565/2803" severity error;
    assert SOR = '1' report "Error in test case #2565/2803" severity error;
    assert SOL = '1' report "Error in test case #2565/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2566/2803" severity error;
    assert SOR = '1' report "Error in test case #2566/2803" severity error;
    assert SOL = '1' report "Error in test case #2566/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2567/2803" severity error;
    assert SOR = '1' report "Error in test case #2567/2803" severity error;
    assert SOL = '1' report "Error in test case #2567/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2568/2803" severity error;
    assert SOR = '1' report "Error in test case #2568/2803" severity error;
    assert SOL = '1' report "Error in test case #2568/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2569/2803" severity error;
    assert SOR = '1' report "Error in test case #2569/2803" severity error;
    assert SOL = '1' report "Error in test case #2569/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2570/2803" severity error;
    assert SOR = '1' report "Error in test case #2570/2803" severity error;
    assert SOL = '1' report "Error in test case #2570/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2571/2803" severity error;
    assert SOR = '1' report "Error in test case #2571/2803" severity error;
    assert SOL = '1' report "Error in test case #2571/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2572/2803" severity error;
    assert SOR = '1' report "Error in test case #2572/2803" severity error;
    assert SOL = '1' report "Error in test case #2572/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2573/2803" severity error;
    assert SOR = '1' report "Error in test case #2573/2803" severity error;
    assert SOL = '1' report "Error in test case #2573/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2574/2803" severity error;
    assert SOR = '1' report "Error in test case #2574/2803" severity error;
    assert SOL = '1' report "Error in test case #2574/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2575/2803" severity error;
    assert SOR = '1' report "Error in test case #2575/2803" severity error;
    assert SOL = '1' report "Error in test case #2575/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2576/2803" severity error;
    assert SOR = '1' report "Error in test case #2576/2803" severity error;
    assert SOL = '1' report "Error in test case #2576/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2577/2803" severity error;
    assert SOR = '1' report "Error in test case #2577/2803" severity error;
    assert SOL = '1' report "Error in test case #2577/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2578/2803" severity error;
    assert SOR = '1' report "Error in test case #2578/2803" severity error;
    assert SOL = '1' report "Error in test case #2578/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2579/2803" severity error;
    assert SOR = '1' report "Error in test case #2579/2803" severity error;
    assert SOL = '1' report "Error in test case #2579/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2580/2803" severity error;
    assert SOR = '1' report "Error in test case #2580/2803" severity error;
    assert SOL = '1' report "Error in test case #2580/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2581/2803" severity error;
    assert SOR = '1' report "Error in test case #2581/2803" severity error;
    assert SOL = '1' report "Error in test case #2581/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2582/2803" severity error;
    assert SOR = '1' report "Error in test case #2582/2803" severity error;
    assert SOL = '1' report "Error in test case #2582/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2583/2803" severity error;
    assert SOR = '1' report "Error in test case #2583/2803" severity error;
    assert SOL = '1' report "Error in test case #2583/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2584/2803" severity error;
    assert SOR = '1' report "Error in test case #2584/2803" severity error;
    assert SOL = '1' report "Error in test case #2584/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2585/2803" severity error;
    assert SOR = '1' report "Error in test case #2585/2803" severity error;
    assert SOL = '1' report "Error in test case #2585/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2586/2803" severity error;
    assert SOR = '1' report "Error in test case #2586/2803" severity error;
    assert SOL = '1' report "Error in test case #2586/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2587/2803" severity error;
    assert SOR = '1' report "Error in test case #2587/2803" severity error;
    assert SOL = '1' report "Error in test case #2587/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2588/2803" severity error;
    assert SOR = '1' report "Error in test case #2588/2803" severity error;
    assert SOL = '1' report "Error in test case #2588/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2589/2803" severity error;
    assert SOR = '1' report "Error in test case #2589/2803" severity error;
    assert SOL = '1' report "Error in test case #2589/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2590/2803" severity error;
    assert SOR = '1' report "Error in test case #2590/2803" severity error;
    assert SOL = '1' report "Error in test case #2590/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2591/2803" severity error;
    assert SOR = '1' report "Error in test case #2591/2803" severity error;
    assert SOL = '1' report "Error in test case #2591/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2592/2803" severity error;
    assert SOR = '1' report "Error in test case #2592/2803" severity error;
    assert SOL = '1' report "Error in test case #2592/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2593/2803" severity error;
    assert SOR = '1' report "Error in test case #2593/2803" severity error;
    assert SOL = '1' report "Error in test case #2593/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2594/2803" severity error;
    assert SOR = '1' report "Error in test case #2594/2803" severity error;
    assert SOL = '1' report "Error in test case #2594/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2595/2803" severity error;
    assert SOR = '1' report "Error in test case #2595/2803" severity error;
    assert SOL = '1' report "Error in test case #2595/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2596/2803" severity error;
    assert SOR = '1' report "Error in test case #2596/2803" severity error;
    assert SOL = '1' report "Error in test case #2596/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2597/2803" severity error;
    assert SOR = '1' report "Error in test case #2597/2803" severity error;
    assert SOL = '1' report "Error in test case #2597/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2598/2803" severity error;
    assert SOR = '1' report "Error in test case #2598/2803" severity error;
    assert SOL = '1' report "Error in test case #2598/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2599/2803" severity error;
    assert SOR = '1' report "Error in test case #2599/2803" severity error;
    assert SOL = '1' report "Error in test case #2599/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2600/2803" severity error;
    assert SOR = '1' report "Error in test case #2600/2803" severity error;
    assert SOL = '1' report "Error in test case #2600/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2601/2803" severity error;
    assert SOR = '1' report "Error in test case #2601/2803" severity error;
    assert SOL = '1' report "Error in test case #2601/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2602/2803" severity error;
    assert SOR = '1' report "Error in test case #2602/2803" severity error;
    assert SOL = '1' report "Error in test case #2602/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2603/2803" severity error;
    assert SOR = '1' report "Error in test case #2603/2803" severity error;
    assert SOL = '1' report "Error in test case #2603/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2604/2803" severity error;
    assert SOR = '1' report "Error in test case #2604/2803" severity error;
    assert SOL = '1' report "Error in test case #2604/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2605/2803" severity error;
    assert SOR = '1' report "Error in test case #2605/2803" severity error;
    assert SOL = '1' report "Error in test case #2605/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2606/2803" severity error;
    assert SOR = '1' report "Error in test case #2606/2803" severity error;
    assert SOL = '1' report "Error in test case #2606/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2607/2803" severity error;
    assert SOR = '1' report "Error in test case #2607/2803" severity error;
    assert SOL = '1' report "Error in test case #2607/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2608/2803" severity error;
    assert SOR = '1' report "Error in test case #2608/2803" severity error;
    assert SOL = '1' report "Error in test case #2608/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2609/2803" severity error;
    assert SOR = '1' report "Error in test case #2609/2803" severity error;
    assert SOL = '1' report "Error in test case #2609/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2610/2803" severity error;
    assert SOR = '1' report "Error in test case #2610/2803" severity error;
    assert SOL = '1' report "Error in test case #2610/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2611/2803" severity error;
    assert SOR = '1' report "Error in test case #2611/2803" severity error;
    assert SOL = '1' report "Error in test case #2611/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2612/2803" severity error;
    assert SOR = '1' report "Error in test case #2612/2803" severity error;
    assert SOL = '1' report "Error in test case #2612/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2613/2803" severity error;
    assert SOR = '1' report "Error in test case #2613/2803" severity error;
    assert SOL = '1' report "Error in test case #2613/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2614/2803" severity error;
    assert SOR = '1' report "Error in test case #2614/2803" severity error;
    assert SOL = '1' report "Error in test case #2614/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2615/2803" severity error;
    assert SOR = '1' report "Error in test case #2615/2803" severity error;
    assert SOL = '1' report "Error in test case #2615/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2616/2803" severity error;
    assert SOR = '1' report "Error in test case #2616/2803" severity error;
    assert SOL = '1' report "Error in test case #2616/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2617/2803" severity error;
    assert SOR = '1' report "Error in test case #2617/2803" severity error;
    assert SOL = '1' report "Error in test case #2617/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2618/2803" severity error;
    assert SOR = '1' report "Error in test case #2618/2803" severity error;
    assert SOL = '1' report "Error in test case #2618/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2619/2803" severity error;
    assert SOR = '1' report "Error in test case #2619/2803" severity error;
    assert SOL = '1' report "Error in test case #2619/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2620/2803" severity error;
    assert SOR = '1' report "Error in test case #2620/2803" severity error;
    assert SOL = '1' report "Error in test case #2620/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2621/2803" severity error;
    assert SOR = '1' report "Error in test case #2621/2803" severity error;
    assert SOL = '1' report "Error in test case #2621/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2622/2803" severity error;
    assert SOR = '1' report "Error in test case #2622/2803" severity error;
    assert SOL = '1' report "Error in test case #2622/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2623/2803" severity error;
    assert SOR = '1' report "Error in test case #2623/2803" severity error;
    assert SOL = '1' report "Error in test case #2623/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2624/2803" severity error;
    assert SOR = '1' report "Error in test case #2624/2803" severity error;
    assert SOL = '1' report "Error in test case #2624/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2625/2803" severity error;
    assert SOR = '1' report "Error in test case #2625/2803" severity error;
    assert SOL = '1' report "Error in test case #2625/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2626/2803" severity error;
    assert SOR = '1' report "Error in test case #2626/2803" severity error;
    assert SOL = '1' report "Error in test case #2626/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2627/2803" severity error;
    assert SOR = '1' report "Error in test case #2627/2803" severity error;
    assert SOL = '1' report "Error in test case #2627/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2628/2803" severity error;
    assert SOR = '1' report "Error in test case #2628/2803" severity error;
    assert SOL = '1' report "Error in test case #2628/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2629/2803" severity error;
    assert SOR = '1' report "Error in test case #2629/2803" severity error;
    assert SOL = '1' report "Error in test case #2629/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2630/2803" severity error;
    assert SOR = '1' report "Error in test case #2630/2803" severity error;
    assert SOL = '1' report "Error in test case #2630/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2631/2803" severity error;
    assert SOR = '1' report "Error in test case #2631/2803" severity error;
    assert SOL = '1' report "Error in test case #2631/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2632/2803" severity error;
    assert SOR = '1' report "Error in test case #2632/2803" severity error;
    assert SOL = '1' report "Error in test case #2632/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2633/2803" severity error;
    assert SOR = '1' report "Error in test case #2633/2803" severity error;
    assert SOL = '1' report "Error in test case #2633/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2634/2803" severity error;
    assert SOR = '1' report "Error in test case #2634/2803" severity error;
    assert SOL = '1' report "Error in test case #2634/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2635/2803" severity error;
    assert SOR = '1' report "Error in test case #2635/2803" severity error;
    assert SOL = '1' report "Error in test case #2635/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2636/2803" severity error;
    assert SOR = '1' report "Error in test case #2636/2803" severity error;
    assert SOL = '1' report "Error in test case #2636/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2637/2803" severity error;
    assert SOR = '1' report "Error in test case #2637/2803" severity error;
    assert SOL = '1' report "Error in test case #2637/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2638/2803" severity error;
    assert SOR = '1' report "Error in test case #2638/2803" severity error;
    assert SOL = '1' report "Error in test case #2638/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2639/2803" severity error;
    assert SOR = '1' report "Error in test case #2639/2803" severity error;
    assert SOL = '1' report "Error in test case #2639/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2640/2803" severity error;
    assert SOR = '1' report "Error in test case #2640/2803" severity error;
    assert SOL = '1' report "Error in test case #2640/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2641/2803" severity error;
    assert SOR = '1' report "Error in test case #2641/2803" severity error;
    assert SOL = '1' report "Error in test case #2641/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2642/2803" severity error;
    assert SOR = '1' report "Error in test case #2642/2803" severity error;
    assert SOL = '1' report "Error in test case #2642/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2643/2803" severity error;
    assert SOR = '1' report "Error in test case #2643/2803" severity error;
    assert SOL = '1' report "Error in test case #2643/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2644/2803" severity error;
    assert SOR = '1' report "Error in test case #2644/2803" severity error;
    assert SOL = '1' report "Error in test case #2644/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2645/2803" severity error;
    assert SOR = '1' report "Error in test case #2645/2803" severity error;
    assert SOL = '1' report "Error in test case #2645/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2646/2803" severity error;
    assert SOR = '1' report "Error in test case #2646/2803" severity error;
    assert SOL = '1' report "Error in test case #2646/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2647/2803" severity error;
    assert SOR = '1' report "Error in test case #2647/2803" severity error;
    assert SOL = '1' report "Error in test case #2647/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2648/2803" severity error;
    assert SOR = '1' report "Error in test case #2648/2803" severity error;
    assert SOL = '1' report "Error in test case #2648/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2649/2803" severity error;
    assert SOR = '1' report "Error in test case #2649/2803" severity error;
    assert SOL = '1' report "Error in test case #2649/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2650/2803" severity error;
    assert SOR = '1' report "Error in test case #2650/2803" severity error;
    assert SOL = '1' report "Error in test case #2650/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2651/2803" severity error;
    assert SOR = '1' report "Error in test case #2651/2803" severity error;
    assert SOL = '1' report "Error in test case #2651/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2652/2803" severity error;
    assert SOR = '1' report "Error in test case #2652/2803" severity error;
    assert SOL = '1' report "Error in test case #2652/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2653/2803" severity error;
    assert SOR = '1' report "Error in test case #2653/2803" severity error;
    assert SOL = '1' report "Error in test case #2653/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2654/2803" severity error;
    assert SOR = '1' report "Error in test case #2654/2803" severity error;
    assert SOL = '1' report "Error in test case #2654/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2655/2803" severity error;
    assert SOR = '1' report "Error in test case #2655/2803" severity error;
    assert SOL = '1' report "Error in test case #2655/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2656/2803" severity error;
    assert SOR = '1' report "Error in test case #2656/2803" severity error;
    assert SOL = '1' report "Error in test case #2656/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2657/2803" severity error;
    assert SOR = '1' report "Error in test case #2657/2803" severity error;
    assert SOL = '1' report "Error in test case #2657/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2658/2803" severity error;
    assert SOR = '1' report "Error in test case #2658/2803" severity error;
    assert SOL = '1' report "Error in test case #2658/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2659/2803" severity error;
    assert SOR = '1' report "Error in test case #2659/2803" severity error;
    assert SOL = '1' report "Error in test case #2659/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2660/2803" severity error;
    assert SOR = '1' report "Error in test case #2660/2803" severity error;
    assert SOL = '1' report "Error in test case #2660/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2661/2803" severity error;
    assert SOR = '1' report "Error in test case #2661/2803" severity error;
    assert SOL = '1' report "Error in test case #2661/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2662/2803" severity error;
    assert SOR = '1' report "Error in test case #2662/2803" severity error;
    assert SOL = '1' report "Error in test case #2662/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2663/2803" severity error;
    assert SOR = '1' report "Error in test case #2663/2803" severity error;
    assert SOL = '1' report "Error in test case #2663/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2664/2803" severity error;
    assert SOR = '1' report "Error in test case #2664/2803" severity error;
    assert SOL = '1' report "Error in test case #2664/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2665/2803" severity error;
    assert SOR = '1' report "Error in test case #2665/2803" severity error;
    assert SOL = '1' report "Error in test case #2665/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2666/2803" severity error;
    assert SOR = '1' report "Error in test case #2666/2803" severity error;
    assert SOL = '1' report "Error in test case #2666/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2667/2803" severity error;
    assert SOR = '1' report "Error in test case #2667/2803" severity error;
    assert SOL = '1' report "Error in test case #2667/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2668/2803" severity error;
    assert SOR = '1' report "Error in test case #2668/2803" severity error;
    assert SOL = '1' report "Error in test case #2668/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2669/2803" severity error;
    assert SOR = '1' report "Error in test case #2669/2803" severity error;
    assert SOL = '1' report "Error in test case #2669/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2670/2803" severity error;
    assert SOR = '1' report "Error in test case #2670/2803" severity error;
    assert SOL = '1' report "Error in test case #2670/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2671/2803" severity error;
    assert SOR = '1' report "Error in test case #2671/2803" severity error;
    assert SOL = '1' report "Error in test case #2671/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2672/2803" severity error;
    assert SOR = '1' report "Error in test case #2672/2803" severity error;
    assert SOL = '1' report "Error in test case #2672/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2673/2803" severity error;
    assert SOR = '1' report "Error in test case #2673/2803" severity error;
    assert SOL = '1' report "Error in test case #2673/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2674/2803" severity error;
    assert SOR = '1' report "Error in test case #2674/2803" severity error;
    assert SOL = '1' report "Error in test case #2674/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2675/2803" severity error;
    assert SOR = '1' report "Error in test case #2675/2803" severity error;
    assert SOL = '1' report "Error in test case #2675/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2676/2803" severity error;
    assert SOR = '1' report "Error in test case #2676/2803" severity error;
    assert SOL = '1' report "Error in test case #2676/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2677/2803" severity error;
    assert SOR = '1' report "Error in test case #2677/2803" severity error;
    assert SOL = '1' report "Error in test case #2677/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2678/2803" severity error;
    assert SOR = '1' report "Error in test case #2678/2803" severity error;
    assert SOL = '1' report "Error in test case #2678/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2679/2803" severity error;
    assert SOR = '0' report "Error in test case #2679/2803" severity error;
    assert SOL = '0' report "Error in test case #2679/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2680/2803" severity error;
    assert SOR = '0' report "Error in test case #2680/2803" severity error;
    assert SOL = '0' report "Error in test case #2680/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2681/2803" severity error;
    assert SOR = '0' report "Error in test case #2681/2803" severity error;
    assert SOL = '0' report "Error in test case #2681/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2682/2803" severity error;
    assert SOR = '0' report "Error in test case #2682/2803" severity error;
    assert SOL = '0' report "Error in test case #2682/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2683/2803" severity error;
    assert SOR = '0' report "Error in test case #2683/2803" severity error;
    assert SOL = '0' report "Error in test case #2683/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2684/2803" severity error;
    assert SOR = '0' report "Error in test case #2684/2803" severity error;
    assert SOL = '0' report "Error in test case #2684/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2685/2803" severity error;
    assert SOR = '0' report "Error in test case #2685/2803" severity error;
    assert SOL = '0' report "Error in test case #2685/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2686/2803" severity error;
    assert SOR = '0' report "Error in test case #2686/2803" severity error;
    assert SOL = '0' report "Error in test case #2686/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2687/2803" severity error;
    assert SOR = '0' report "Error in test case #2687/2803" severity error;
    assert SOL = '0' report "Error in test case #2687/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2688/2803" severity error;
    assert SOR = '0' report "Error in test case #2688/2803" severity error;
    assert SOL = '0' report "Error in test case #2688/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2689/2803" severity error;
    assert SOR = '0' report "Error in test case #2689/2803" severity error;
    assert SOL = '0' report "Error in test case #2689/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2690/2803" severity error;
    assert SOR = '0' report "Error in test case #2690/2803" severity error;
    assert SOL = '0' report "Error in test case #2690/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2691/2803" severity error;
    assert SOR = '0' report "Error in test case #2691/2803" severity error;
    assert SOL = '0' report "Error in test case #2691/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2692/2803" severity error;
    assert SOR = '0' report "Error in test case #2692/2803" severity error;
    assert SOL = '0' report "Error in test case #2692/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2693/2803" severity error;
    assert SOR = '0' report "Error in test case #2693/2803" severity error;
    assert SOL = '0' report "Error in test case #2693/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2694/2803" severity error;
    assert SOR = '0' report "Error in test case #2694/2803" severity error;
    assert SOL = '0' report "Error in test case #2694/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2695/2803" severity error;
    assert SOR = '0' report "Error in test case #2695/2803" severity error;
    assert SOL = '0' report "Error in test case #2695/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2696/2803" severity error;
    assert SOR = '0' report "Error in test case #2696/2803" severity error;
    assert SOL = '0' report "Error in test case #2696/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2697/2803" severity error;
    assert SOR = '1' report "Error in test case #2697/2803" severity error;
    assert SOL = '1' report "Error in test case #2697/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2698/2803" severity error;
    assert SOR = '1' report "Error in test case #2698/2803" severity error;
    assert SOL = '1' report "Error in test case #2698/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2699/2803" severity error;
    assert SOR = '1' report "Error in test case #2699/2803" severity error;
    assert SOL = '1' report "Error in test case #2699/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2700/2803" severity error;
    assert SOR = '1' report "Error in test case #2700/2803" severity error;
    assert SOL = '1' report "Error in test case #2700/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2701/2803" severity error;
    assert SOR = '1' report "Error in test case #2701/2803" severity error;
    assert SOL = '1' report "Error in test case #2701/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2702/2803" severity error;
    assert SOR = '1' report "Error in test case #2702/2803" severity error;
    assert SOL = '1' report "Error in test case #2702/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2703/2803" severity error;
    assert SOR = '1' report "Error in test case #2703/2803" severity error;
    assert SOL = '1' report "Error in test case #2703/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2704/2803" severity error;
    assert SOR = '1' report "Error in test case #2704/2803" severity error;
    assert SOL = '1' report "Error in test case #2704/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2705/2803" severity error;
    assert SOR = '1' report "Error in test case #2705/2803" severity error;
    assert SOL = '1' report "Error in test case #2705/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2706/2803" severity error;
    assert SOR = '1' report "Error in test case #2706/2803" severity error;
    assert SOL = '1' report "Error in test case #2706/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2707/2803" severity error;
    assert SOR = '1' report "Error in test case #2707/2803" severity error;
    assert SOL = '1' report "Error in test case #2707/2803" severity error;

    CLK <= '0';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2708/2803" severity error;
    assert SOR = '0' report "Error in test case #2708/2803" severity error;
    assert SOL = '0' report "Error in test case #2708/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2709/2803" severity error;
    assert SOR = '0' report "Error in test case #2709/2803" severity error;
    assert SOL = '0' report "Error in test case #2709/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2710/2803" severity error;
    assert SOR = '0' report "Error in test case #2710/2803" severity error;
    assert SOL = '0' report "Error in test case #2710/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2711/2803" severity error;
    assert SOR = '0' report "Error in test case #2711/2803" severity error;
    assert SOL = '0' report "Error in test case #2711/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2712/2803" severity error;
    assert SOR = '0' report "Error in test case #2712/2803" severity error;
    assert SOL = '0' report "Error in test case #2712/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2713/2803" severity error;
    assert SOR = '0' report "Error in test case #2713/2803" severity error;
    assert SOL = '0' report "Error in test case #2713/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2714/2803" severity error;
    assert SOR = '0' report "Error in test case #2714/2803" severity error;
    assert SOL = '0' report "Error in test case #2714/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2715/2803" severity error;
    assert SOR = '0' report "Error in test case #2715/2803" severity error;
    assert SOL = '0' report "Error in test case #2715/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2716/2803" severity error;
    assert SOR = '0' report "Error in test case #2716/2803" severity error;
    assert SOL = '0' report "Error in test case #2716/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2717/2803" severity error;
    assert SOR = '0' report "Error in test case #2717/2803" severity error;
    assert SOL = '0' report "Error in test case #2717/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2718/2803" severity error;
    assert SOR = '0' report "Error in test case #2718/2803" severity error;
    assert SOL = '0' report "Error in test case #2718/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2719/2803" severity error;
    assert SOR = '0' report "Error in test case #2719/2803" severity error;
    assert SOL = '0' report "Error in test case #2719/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2720/2803" severity error;
    assert SOR = '0' report "Error in test case #2720/2803" severity error;
    assert SOL = '0' report "Error in test case #2720/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2721/2803" severity error;
    assert SOR = '0' report "Error in test case #2721/2803" severity error;
    assert SOL = '0' report "Error in test case #2721/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2722/2803" severity error;
    assert SOR = '0' report "Error in test case #2722/2803" severity error;
    assert SOL = '0' report "Error in test case #2722/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2723/2803" severity error;
    assert SOR = '0' report "Error in test case #2723/2803" severity error;
    assert SOL = '0' report "Error in test case #2723/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2724/2803" severity error;
    assert SOR = '0' report "Error in test case #2724/2803" severity error;
    assert SOL = '0' report "Error in test case #2724/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2725/2803" severity error;
    assert SOR = '0' report "Error in test case #2725/2803" severity error;
    assert SOL = '0' report "Error in test case #2725/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2726/2803" severity error;
    assert SOR = '0' report "Error in test case #2726/2803" severity error;
    assert SOL = '0' report "Error in test case #2726/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2727/2803" severity error;
    assert SOR = '0' report "Error in test case #2727/2803" severity error;
    assert SOL = '0' report "Error in test case #2727/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2728/2803" severity error;
    assert SOR = '0' report "Error in test case #2728/2803" severity error;
    assert SOL = '0' report "Error in test case #2728/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2729/2803" severity error;
    assert SOR = '0' report "Error in test case #2729/2803" severity error;
    assert SOL = '0' report "Error in test case #2729/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2730/2803" severity error;
    assert SOR = '0' report "Error in test case #2730/2803" severity error;
    assert SOL = '0' report "Error in test case #2730/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2731/2803" severity error;
    assert SOR = '0' report "Error in test case #2731/2803" severity error;
    assert SOL = '0' report "Error in test case #2731/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2732/2803" severity error;
    assert SOR = '0' report "Error in test case #2732/2803" severity error;
    assert SOL = '0' report "Error in test case #2732/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2733/2803" severity error;
    assert SOR = '0' report "Error in test case #2733/2803" severity error;
    assert SOL = '0' report "Error in test case #2733/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2734/2803" severity error;
    assert SOR = '0' report "Error in test case #2734/2803" severity error;
    assert SOL = '0' report "Error in test case #2734/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2735/2803" severity error;
    assert SOR = '0' report "Error in test case #2735/2803" severity error;
    assert SOL = '0' report "Error in test case #2735/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2736/2803" severity error;
    assert SOR = '0' report "Error in test case #2736/2803" severity error;
    assert SOL = '0' report "Error in test case #2736/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2737/2803" severity error;
    assert SOR = '0' report "Error in test case #2737/2803" severity error;
    assert SOL = '0' report "Error in test case #2737/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2738/2803" severity error;
    assert SOR = '0' report "Error in test case #2738/2803" severity error;
    assert SOL = '0' report "Error in test case #2738/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2739/2803" severity error;
    assert SOR = '0' report "Error in test case #2739/2803" severity error;
    assert SOL = '0' report "Error in test case #2739/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2740/2803" severity error;
    assert SOR = '0' report "Error in test case #2740/2803" severity error;
    assert SOL = '0' report "Error in test case #2740/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000101";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2741/2803" severity error;
    assert SOR = '0' report "Error in test case #2741/2803" severity error;
    assert SOL = '0' report "Error in test case #2741/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2742/2803" severity error;
    assert SOR = '0' report "Error in test case #2742/2803" severity error;
    assert SOL = '0' report "Error in test case #2742/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2743/2803" severity error;
    assert SOR = '0' report "Error in test case #2743/2803" severity error;
    assert SOL = '0' report "Error in test case #2743/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2744/2803" severity error;
    assert SOR = '0' report "Error in test case #2744/2803" severity error;
    assert SOL = '0' report "Error in test case #2744/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2745/2803" severity error;
    assert SOR = '0' report "Error in test case #2745/2803" severity error;
    assert SOL = '0' report "Error in test case #2745/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2746/2803" severity error;
    assert SOR = '0' report "Error in test case #2746/2803" severity error;
    assert SOL = '0' report "Error in test case #2746/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2747/2803" severity error;
    assert SOR = '0' report "Error in test case #2747/2803" severity error;
    assert SOL = '0' report "Error in test case #2747/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2748/2803" severity error;
    assert SOR = '0' report "Error in test case #2748/2803" severity error;
    assert SOL = '0' report "Error in test case #2748/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2749/2803" severity error;
    assert SOR = '0' report "Error in test case #2749/2803" severity error;
    assert SOL = '0' report "Error in test case #2749/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2750/2803" severity error;
    assert SOR = '0' report "Error in test case #2750/2803" severity error;
    assert SOL = '0' report "Error in test case #2750/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2751/2803" severity error;
    assert SOR = '0' report "Error in test case #2751/2803" severity error;
    assert SOL = '0' report "Error in test case #2751/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2752/2803" severity error;
    assert SOR = '0' report "Error in test case #2752/2803" severity error;
    assert SOL = '0' report "Error in test case #2752/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2753/2803" severity error;
    assert SOR = '0' report "Error in test case #2753/2803" severity error;
    assert SOL = '0' report "Error in test case #2753/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2754/2803" severity error;
    assert SOR = '1' report "Error in test case #2754/2803" severity error;
    assert SOL = '1' report "Error in test case #2754/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2755/2803" severity error;
    assert SOR = '1' report "Error in test case #2755/2803" severity error;
    assert SOL = '1' report "Error in test case #2755/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2756/2803" severity error;
    assert SOR = '1' report "Error in test case #2756/2803" severity error;
    assert SOL = '1' report "Error in test case #2756/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2757/2803" severity error;
    assert SOR = '1' report "Error in test case #2757/2803" severity error;
    assert SOL = '1' report "Error in test case #2757/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2758/2803" severity error;
    assert SOR = '1' report "Error in test case #2758/2803" severity error;
    assert SOL = '1' report "Error in test case #2758/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2759/2803" severity error;
    assert SOR = '1' report "Error in test case #2759/2803" severity error;
    assert SOL = '1' report "Error in test case #2759/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2760/2803" severity error;
    assert SOR = '1' report "Error in test case #2760/2803" severity error;
    assert SOL = '1' report "Error in test case #2760/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2761/2803" severity error;
    assert SOR = '1' report "Error in test case #2761/2803" severity error;
    assert SOL = '1' report "Error in test case #2761/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '0';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2762/2803" severity error;
    assert SOR = '1' report "Error in test case #2762/2803" severity error;
    assert SOL = '1' report "Error in test case #2762/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2763/2803" severity error;
    assert SOR = '1' report "Error in test case #2763/2803" severity error;
    assert SOL = '1' report "Error in test case #2763/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2764/2803" severity error;
    assert SOR = '1' report "Error in test case #2764/2803" severity error;
    assert SOL = '1' report "Error in test case #2764/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2765/2803" severity error;
    assert SOR = '1' report "Error in test case #2765/2803" severity error;
    assert SOL = '1' report "Error in test case #2765/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2766/2803" severity error;
    assert SOR = '1' report "Error in test case #2766/2803" severity error;
    assert SOL = '1' report "Error in test case #2766/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2767/2803" severity error;
    assert SOR = '1' report "Error in test case #2767/2803" severity error;
    assert SOL = '1' report "Error in test case #2767/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2768/2803" severity error;
    assert SOR = '1' report "Error in test case #2768/2803" severity error;
    assert SOL = '1' report "Error in test case #2768/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2769/2803" severity error;
    assert SOR = '1' report "Error in test case #2769/2803" severity error;
    assert SOL = '1' report "Error in test case #2769/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2770/2803" severity error;
    assert SOR = '1' report "Error in test case #2770/2803" severity error;
    assert SOL = '1' report "Error in test case #2770/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2771/2803" severity error;
    assert SOR = '1' report "Error in test case #2771/2803" severity error;
    assert SOL = '1' report "Error in test case #2771/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2772/2803" severity error;
    assert SOR = '1' report "Error in test case #2772/2803" severity error;
    assert SOL = '1' report "Error in test case #2772/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2773/2803" severity error;
    assert SOR = '1' report "Error in test case #2773/2803" severity error;
    assert SOL = '1' report "Error in test case #2773/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2774/2803" severity error;
    assert SOR = '1' report "Error in test case #2774/2803" severity error;
    assert SOL = '1' report "Error in test case #2774/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2775/2803" severity error;
    assert SOR = '1' report "Error in test case #2775/2803" severity error;
    assert SOL = '1' report "Error in test case #2775/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "11111111" report "Error in test case #2776/2803" severity error;
    assert SOR = '1' report "Error in test case #2776/2803" severity error;
    assert SOL = '1' report "Error in test case #2776/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2777/2803" severity error;
    assert SOR = '0' report "Error in test case #2777/2803" severity error;
    assert SOL = '0' report "Error in test case #2777/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2778/2803" severity error;
    assert SOR = '0' report "Error in test case #2778/2803" severity error;
    assert SOL = '0' report "Error in test case #2778/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2779/2803" severity error;
    assert SOR = '0' report "Error in test case #2779/2803" severity error;
    assert SOL = '0' report "Error in test case #2779/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2780/2803" severity error;
    assert SOR = '0' report "Error in test case #2780/2803" severity error;
    assert SOL = '0' report "Error in test case #2780/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2781/2803" severity error;
    assert SOR = '0' report "Error in test case #2781/2803" severity error;
    assert SOL = '0' report "Error in test case #2781/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2782/2803" severity error;
    assert SOR = '0' report "Error in test case #2782/2803" severity error;
    assert SOL = '0' report "Error in test case #2782/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2783/2803" severity error;
    assert SOR = '0' report "Error in test case #2783/2803" severity error;
    assert SOL = '0' report "Error in test case #2783/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2784/2803" severity error;
    assert SOR = '0' report "Error in test case #2784/2803" severity error;
    assert SOL = '0' report "Error in test case #2784/2803" severity error;

    CLK <= '1';
    RSTn <= '0';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2785/2803" severity error;
    assert SOR = '0' report "Error in test case #2785/2803" severity error;
    assert SOL = '0' report "Error in test case #2785/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2786/2803" severity error;
    assert SOR = '0' report "Error in test case #2786/2803" severity error;
    assert SOL = '0' report "Error in test case #2786/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2787/2803" severity error;
    assert SOR = '0' report "Error in test case #2787/2803" severity error;
    assert SOL = '0' report "Error in test case #2787/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000101";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2788/2803" severity error;
    assert SOR = '0' report "Error in test case #2788/2803" severity error;
    assert SOL = '0' report "Error in test case #2788/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000000";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2789/2803" severity error;
    assert SOR = '0' report "Error in test case #2789/2803" severity error;
    assert SOL = '0' report "Error in test case #2789/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2790/2803" severity error;
    assert SOR = '0' report "Error in test case #2790/2803" severity error;
    assert SOL = '0' report "Error in test case #2790/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2791/2803" severity error;
    assert SOR = '0' report "Error in test case #2791/2803" severity error;
    assert SOL = '0' report "Error in test case #2791/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2792/2803" severity error;
    assert SOR = '0' report "Error in test case #2792/2803" severity error;
    assert SOL = '0' report "Error in test case #2792/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000110";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2793/2803" severity error;
    assert SOR = '0' report "Error in test case #2793/2803" severity error;
    assert SOL = '0' report "Error in test case #2793/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000001";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2794/2803" severity error;
    assert SOR = '0' report "Error in test case #2794/2803" severity error;
    assert SOL = '0' report "Error in test case #2794/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2795/2803" severity error;
    assert SOR = '0' report "Error in test case #2795/2803" severity error;
    assert SOL = '0' report "Error in test case #2795/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000100";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2796/2803" severity error;
    assert SOR = '0' report "Error in test case #2796/2803" severity error;
    assert SOL = '0' report "Error in test case #2796/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000000";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2797/2803" severity error;
    assert SOR = '0' report "Error in test case #2797/2803" severity error;
    assert SOL = '0' report "Error in test case #2797/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '0';
    Pi <= "00000010";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2798/2803" severity error;
    assert SOR = '0' report "Error in test case #2798/2803" severity error;
    assert SOL = '0' report "Error in test case #2798/2803" severity error;

    CLK <= '0';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2799/2803" severity error;
    assert SOR = '0' report "Error in test case #2799/2803" severity error;
    assert SOL = '0' report "Error in test case #2799/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000110";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2800/2803" severity error;
    assert SOR = '0' report "Error in test case #2800/2803" severity error;
    assert SOL = '0' report "Error in test case #2800/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2801/2803" severity error;
    assert SOR = '0' report "Error in test case #2801/2803" severity error;
    assert SOL = '0' report "Error in test case #2801/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000011";
    SSL <= '1';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2802/2803" severity error;
    assert SOR = '0' report "Error in test case #2802/2803" severity error;
    assert SOL = '0' report "Error in test case #2802/2803" severity error;

    CLK <= '1';
    RSTn <= '1';
    SETn <= '1';
    SEL <= "110";
    SSR <= '1';
    Pi <= "00000111";
    SSL <= '0';
    wait for 10 ns;
    assert Qo = "00000000" report "Error in test case #2803/2803" severity error;
    assert SOR = '0' report "Error in test case #2803/2803" severity error;
    assert SOL = '0' report "Error in test case #2803/2803" severity error;

    wait;
end process;
	
END universal_register_arch;